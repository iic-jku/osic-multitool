magic
tech sky130A
magscale 1 2
timestamp 1640642158
<< viali >>
rect 1501 8585 1535 8619
rect 4905 8585 4939 8619
rect 1685 8449 1719 8483
rect 4721 8449 4755 8483
rect 4629 7361 4663 7395
rect 4537 7157 4571 7191
rect 2145 6817 2179 6851
rect 2237 6749 2271 6783
rect 3985 6749 4019 6783
rect 4813 6681 4847 6715
rect 3893 6613 3927 6647
rect 4721 6613 4755 6647
rect 4997 6409 5031 6443
rect 3902 6341 3936 6375
rect 2145 6273 2179 6307
rect 2237 6273 2271 6307
rect 4629 6273 4663 6307
rect 4721 6273 4755 6307
rect 4169 6205 4203 6239
rect 2789 6069 2823 6103
rect 4629 6069 4663 6103
rect 3249 5729 3283 5763
rect 4261 5729 4295 5763
rect 3985 5661 4019 5695
rect 4169 5661 4203 5695
rect 4353 5661 4387 5695
rect 4537 5661 4571 5695
rect 3004 5593 3038 5627
rect 3801 5593 3835 5627
rect 1869 5525 1903 5559
rect 2973 5253 3007 5287
rect 2237 5185 2271 5219
rect 2513 5117 2547 5151
rect 2053 4981 2087 5015
rect 2421 4981 2455 5015
rect 4261 4981 4295 5015
rect 1593 4777 1627 4811
rect 3801 4777 3835 4811
rect 4169 4641 4203 4675
rect 2973 4573 3007 4607
rect 3985 4573 4019 4607
rect 4261 4573 4295 4607
rect 4353 4573 4387 4607
rect 4537 4573 4571 4607
rect 2706 4505 2740 4539
rect 2053 4233 2087 4267
rect 2053 4097 2087 4131
rect 2329 4097 2363 4131
rect 3065 4097 3099 4131
rect 3157 4097 3191 4131
rect 3884 4097 3918 4131
rect 3617 4029 3651 4063
rect 2145 3961 2179 3995
rect 4997 3893 5031 3927
rect 2421 3689 2455 3723
rect 3893 3689 3927 3723
rect 4445 3689 4479 3723
rect 2513 3485 2547 3519
rect 3985 3485 4019 3519
rect 4445 3485 4479 3519
rect 4629 3485 4663 3519
rect 4813 3145 4847 3179
rect 4997 3009 5031 3043
rect 1685 2397 1719 2431
rect 4721 2397 4755 2431
rect 1501 2261 1535 2295
rect 4905 2261 4939 2295
<< metal1 >>
rect 1104 8730 5704 8752
rect 1104 8678 2491 8730
rect 2543 8678 2555 8730
rect 2607 8678 2619 8730
rect 2671 8678 2683 8730
rect 2735 8678 2747 8730
rect 2799 8678 4033 8730
rect 4085 8678 4097 8730
rect 4149 8678 4161 8730
rect 4213 8678 4225 8730
rect 4277 8678 4289 8730
rect 4341 8678 5704 8730
rect 1104 8656 5704 8678
rect 658 8576 664 8628
rect 716 8616 722 8628
rect 1489 8619 1547 8625
rect 1489 8616 1501 8619
rect 716 8588 1501 8616
rect 716 8576 722 8588
rect 1489 8585 1501 8588
rect 1535 8585 1547 8619
rect 1489 8579 1547 8585
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 6454 8616 6460 8628
rect 4939 8588 6460 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2130 8480 2136 8492
rect 1719 8452 2136 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 4614 8440 4620 8492
rect 4672 8480 4678 8492
rect 4709 8483 4767 8489
rect 4709 8480 4721 8483
rect 4672 8452 4721 8480
rect 4672 8440 4678 8452
rect 4709 8449 4721 8452
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 1104 8186 5704 8208
rect 1104 8134 1721 8186
rect 1773 8134 1785 8186
rect 1837 8134 1849 8186
rect 1901 8134 1913 8186
rect 1965 8134 1977 8186
rect 2029 8134 3262 8186
rect 3314 8134 3326 8186
rect 3378 8134 3390 8186
rect 3442 8134 3454 8186
rect 3506 8134 3518 8186
rect 3570 8134 4804 8186
rect 4856 8134 4868 8186
rect 4920 8134 4932 8186
rect 4984 8134 4996 8186
rect 5048 8134 5060 8186
rect 5112 8134 5704 8186
rect 1104 8112 5704 8134
rect 1104 7642 5704 7664
rect 1104 7590 2491 7642
rect 2543 7590 2555 7642
rect 2607 7590 2619 7642
rect 2671 7590 2683 7642
rect 2735 7590 2747 7642
rect 2799 7590 4033 7642
rect 4085 7590 4097 7642
rect 4149 7590 4161 7642
rect 4213 7590 4225 7642
rect 4277 7590 4289 7642
rect 4341 7590 5704 7642
rect 1104 7568 5704 7590
rect 4614 7392 4620 7404
rect 4575 7364 4620 7392
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 4488 7160 4537 7188
rect 4488 7148 4494 7160
rect 4525 7157 4537 7160
rect 4571 7157 4583 7191
rect 4525 7151 4583 7157
rect 1104 7098 5704 7120
rect 1104 7046 1721 7098
rect 1773 7046 1785 7098
rect 1837 7046 1849 7098
rect 1901 7046 1913 7098
rect 1965 7046 1977 7098
rect 2029 7046 3262 7098
rect 3314 7046 3326 7098
rect 3378 7046 3390 7098
rect 3442 7046 3454 7098
rect 3506 7046 3518 7098
rect 3570 7046 4804 7098
rect 4856 7046 4868 7098
rect 4920 7046 4932 7098
rect 4984 7046 4996 7098
rect 5048 7046 5060 7098
rect 5112 7046 5704 7098
rect 1104 7024 5704 7046
rect 2133 6851 2191 6857
rect 2133 6817 2145 6851
rect 2179 6848 2191 6851
rect 5166 6848 5172 6860
rect 2179 6820 5172 6848
rect 2179 6817 2191 6820
rect 2133 6811 2191 6817
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2314 6780 2320 6792
rect 2271 6752 2320 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 3878 6740 3884 6792
rect 3936 6740 3942 6792
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6780 4031 6783
rect 4614 6780 4620 6792
rect 4019 6752 4620 6780
rect 4019 6749 4031 6752
rect 3973 6743 4031 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 3896 6712 3924 6740
rect 4801 6715 4859 6721
rect 4801 6712 4813 6715
rect 3896 6684 4813 6712
rect 4801 6681 4813 6684
rect 4847 6681 4859 6715
rect 4801 6675 4859 6681
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3752 6616 3893 6644
rect 3752 6604 3758 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 3881 6607 3939 6613
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 4580 6616 4721 6644
rect 4580 6604 4586 6616
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 1104 6554 5704 6576
rect 1104 6502 2491 6554
rect 2543 6502 2555 6554
rect 2607 6502 2619 6554
rect 2671 6502 2683 6554
rect 2735 6502 2747 6554
rect 2799 6502 4033 6554
rect 4085 6502 4097 6554
rect 4149 6502 4161 6554
rect 4213 6502 4225 6554
rect 4277 6502 4289 6554
rect 4341 6502 5704 6554
rect 1104 6480 5704 6502
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 3660 6412 4016 6440
rect 3660 6400 3666 6412
rect 3786 6332 3792 6384
rect 3844 6372 3850 6384
rect 3890 6375 3948 6381
rect 3890 6372 3902 6375
rect 3844 6344 3902 6372
rect 3844 6332 3850 6344
rect 3890 6341 3902 6344
rect 3936 6341 3948 6375
rect 3988 6372 4016 6412
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 4985 6443 5043 6449
rect 4985 6440 4997 6443
rect 4672 6412 4997 6440
rect 4672 6400 4678 6412
rect 4985 6409 4997 6412
rect 5031 6409 5043 6443
rect 4985 6403 5043 6409
rect 3988 6344 4752 6372
rect 3890 6335 3948 6341
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 2130 6304 2136 6316
rect 1636 6276 2136 6304
rect 1636 6264 1642 6276
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 2222 6264 2228 6316
rect 2280 6304 2286 6316
rect 4724 6313 4752 6344
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 2280 6276 4629 6304
rect 2280 6264 2286 6276
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4154 6236 4160 6248
rect 4115 6208 4160 6236
rect 4154 6196 4160 6208
rect 4212 6236 4218 6248
rect 4522 6236 4528 6248
rect 4212 6208 4528 6236
rect 4212 6196 4218 6208
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 2866 6100 2872 6112
rect 2823 6072 2872 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 4580 6072 4629 6100
rect 4580 6060 4586 6072
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 4617 6063 4675 6069
rect 1104 6010 5704 6032
rect 1104 5958 1721 6010
rect 1773 5958 1785 6010
rect 1837 5958 1849 6010
rect 1901 5958 1913 6010
rect 1965 5958 1977 6010
rect 2029 5958 3262 6010
rect 3314 5958 3326 6010
rect 3378 5958 3390 6010
rect 3442 5958 3454 6010
rect 3506 5958 3518 6010
rect 3570 5958 4804 6010
rect 4856 5958 4868 6010
rect 4920 5958 4932 6010
rect 4984 5958 4996 6010
rect 5048 5958 5060 6010
rect 5112 5958 5704 6010
rect 1104 5936 5704 5958
rect 4154 5828 4160 5840
rect 3252 5800 4160 5828
rect 3252 5769 3280 5800
rect 4154 5788 4160 5800
rect 4212 5788 4218 5840
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5729 3295 5763
rect 3694 5760 3700 5772
rect 3237 5723 3295 5729
rect 3436 5732 3700 5760
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3436 5692 3464 5732
rect 3694 5720 3700 5732
rect 3752 5760 3758 5772
rect 4249 5763 4307 5769
rect 3752 5732 4200 5760
rect 3752 5720 3758 5732
rect 4172 5701 4200 5732
rect 4249 5729 4261 5763
rect 4295 5760 4307 5763
rect 4614 5760 4620 5772
rect 4295 5732 4620 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 3200 5664 3464 5692
rect 3973 5695 4031 5701
rect 3200 5652 3206 5664
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 4430 5692 4436 5704
rect 4387 5664 4436 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 2992 5627 3050 5633
rect 2992 5593 3004 5627
rect 3038 5624 3050 5627
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 3038 5596 3801 5624
rect 3038 5593 3050 5596
rect 2992 5587 3050 5593
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 3789 5587 3847 5593
rect 3988 5624 4016 5655
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 5166 5692 5172 5704
rect 4571 5664 5172 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 4706 5624 4712 5636
rect 3988 5596 4712 5624
rect 1857 5559 1915 5565
rect 1857 5525 1869 5559
rect 1903 5556 1915 5559
rect 3988 5556 4016 5596
rect 4706 5584 4712 5596
rect 4764 5584 4770 5636
rect 1903 5528 4016 5556
rect 1903 5525 1915 5528
rect 1857 5519 1915 5525
rect 1104 5466 5704 5488
rect 1104 5414 2491 5466
rect 2543 5414 2555 5466
rect 2607 5414 2619 5466
rect 2671 5414 2683 5466
rect 2735 5414 2747 5466
rect 2799 5414 4033 5466
rect 4085 5414 4097 5466
rect 4149 5414 4161 5466
rect 4213 5414 4225 5466
rect 4277 5414 4289 5466
rect 4341 5414 5704 5466
rect 1104 5392 5704 5414
rect 2958 5284 2964 5296
rect 2919 5256 2964 5284
rect 2958 5244 2964 5256
rect 3016 5244 3022 5296
rect 2222 5216 2228 5228
rect 2183 5188 2228 5216
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 3602 5148 3608 5160
rect 2547 5120 3608 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 2041 5015 2099 5021
rect 2041 4981 2053 5015
rect 2087 5012 2099 5015
rect 2130 5012 2136 5024
rect 2087 4984 2136 5012
rect 2087 4981 2099 4984
rect 2041 4975 2099 4981
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2409 5015 2467 5021
rect 2409 4981 2421 5015
rect 2455 5012 2467 5015
rect 3050 5012 3056 5024
rect 2455 4984 3056 5012
rect 2455 4981 2467 4984
rect 2409 4975 2467 4981
rect 3050 4972 3056 4984
rect 3108 4972 3114 5024
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4249 5015 4307 5021
rect 4249 5012 4261 5015
rect 3936 4984 4261 5012
rect 3936 4972 3942 4984
rect 4249 4981 4261 4984
rect 4295 4981 4307 5015
rect 4249 4975 4307 4981
rect 1104 4922 5704 4944
rect 1104 4870 1721 4922
rect 1773 4870 1785 4922
rect 1837 4870 1849 4922
rect 1901 4870 1913 4922
rect 1965 4870 1977 4922
rect 2029 4870 3262 4922
rect 3314 4870 3326 4922
rect 3378 4870 3390 4922
rect 3442 4870 3454 4922
rect 3506 4870 3518 4922
rect 3570 4870 4804 4922
rect 4856 4870 4868 4922
rect 4920 4870 4932 4922
rect 4984 4870 4996 4922
rect 5048 4870 5060 4922
rect 5112 4870 5704 4922
rect 1104 4848 5704 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4522 4740 4528 4752
rect 4172 4712 4528 4740
rect 3050 4632 3056 4684
rect 3108 4672 3114 4684
rect 4172 4681 4200 4712
rect 4522 4700 4528 4712
rect 4580 4700 4586 4752
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 3108 4644 4169 4672
rect 3108 4632 3114 4644
rect 4157 4641 4169 4644
rect 4203 4641 4215 4675
rect 4157 4635 4215 4641
rect 2958 4604 2964 4616
rect 2919 4576 2964 4604
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 3602 4564 3608 4616
rect 3660 4604 3666 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3660 4576 3985 4604
rect 3660 4564 3666 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4430 4604 4436 4616
rect 4387 4576 4436 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 2038 4496 2044 4548
rect 2096 4536 2102 4548
rect 2694 4539 2752 4545
rect 2694 4536 2706 4539
rect 2096 4508 2706 4536
rect 2096 4496 2102 4508
rect 2694 4505 2706 4508
rect 2740 4505 2752 4539
rect 2694 4499 2752 4505
rect 3694 4496 3700 4548
rect 3752 4536 3758 4548
rect 4264 4536 4292 4567
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4604 4583 4607
rect 5166 4604 5172 4616
rect 4571 4576 5172 4604
rect 4571 4573 4583 4576
rect 4525 4567 4583 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 3752 4508 4292 4536
rect 3752 4496 3758 4508
rect 1104 4378 5704 4400
rect 1104 4326 2491 4378
rect 2543 4326 2555 4378
rect 2607 4326 2619 4378
rect 2671 4326 2683 4378
rect 2735 4326 2747 4378
rect 2799 4326 4033 4378
rect 4085 4326 4097 4378
rect 4149 4326 4161 4378
rect 4213 4326 4225 4378
rect 4277 4326 4289 4378
rect 4341 4326 5704 4378
rect 1104 4304 5704 4326
rect 2038 4264 2044 4276
rect 1999 4236 2044 4264
rect 2038 4224 2044 4236
rect 2096 4224 2102 4276
rect 2884 4168 3188 4196
rect 2884 4140 2912 4168
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2130 4128 2136 4140
rect 2087 4100 2136 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2314 4128 2320 4140
rect 2275 4100 2320 4128
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2866 4088 2872 4140
rect 2924 4088 2930 4140
rect 3050 4128 3056 4140
rect 3011 4100 3056 4128
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 3160 4137 3188 4168
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 3694 4128 3700 4140
rect 3191 4100 3700 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 3872 4131 3930 4137
rect 3872 4097 3884 4131
rect 3918 4128 3930 4131
rect 4430 4128 4436 4140
rect 3918 4100 4436 4128
rect 3918 4097 3930 4100
rect 3872 4091 3930 4097
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 3016 4032 3617 4060
rect 3016 4020 3022 4032
rect 3605 4029 3617 4032
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 2133 3995 2191 4001
rect 2133 3961 2145 3995
rect 2179 3992 2191 3995
rect 3142 3992 3148 4004
rect 2179 3964 3148 3992
rect 2179 3961 2191 3964
rect 2133 3955 2191 3961
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 4985 3927 5043 3933
rect 4985 3924 4997 3927
rect 4580 3896 4997 3924
rect 4580 3884 4586 3896
rect 4985 3893 4997 3896
rect 5031 3893 5043 3927
rect 4985 3887 5043 3893
rect 1104 3834 5704 3856
rect 1104 3782 1721 3834
rect 1773 3782 1785 3834
rect 1837 3782 1849 3834
rect 1901 3782 1913 3834
rect 1965 3782 1977 3834
rect 2029 3782 3262 3834
rect 3314 3782 3326 3834
rect 3378 3782 3390 3834
rect 3442 3782 3454 3834
rect 3506 3782 3518 3834
rect 3570 3782 4804 3834
rect 4856 3782 4868 3834
rect 4920 3782 4932 3834
rect 4984 3782 4996 3834
rect 5048 3782 5060 3834
rect 5112 3782 5704 3834
rect 1104 3760 5704 3782
rect 2409 3723 2467 3729
rect 2409 3689 2421 3723
rect 2455 3720 2467 3723
rect 2958 3720 2964 3732
rect 2455 3692 2964 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 3660 3692 3893 3720
rect 3660 3680 3666 3692
rect 3881 3689 3893 3692
rect 3927 3689 3939 3723
rect 4430 3720 4436 3732
rect 4391 3692 4436 3720
rect 3881 3683 3939 3689
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2372 3556 4660 3584
rect 2372 3544 2378 3556
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 3878 3516 3884 3528
rect 2547 3488 3884 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3516 4031 3519
rect 4430 3516 4436 3528
rect 4019 3488 4436 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 4632 3525 4660 3556
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 4798 3516 4804 3528
rect 4663 3488 4804 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 1104 3290 5704 3312
rect 1104 3238 2491 3290
rect 2543 3238 2555 3290
rect 2607 3238 2619 3290
rect 2671 3238 2683 3290
rect 2735 3238 2747 3290
rect 2799 3238 4033 3290
rect 4085 3238 4097 3290
rect 4149 3238 4161 3290
rect 4213 3238 4225 3290
rect 4277 3238 4289 3290
rect 4341 3238 5704 3290
rect 1104 3216 5704 3238
rect 4798 3176 4804 3188
rect 4759 3148 4804 3176
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3040 5043 3043
rect 5258 3040 5264 3052
rect 5031 3012 5264 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 1104 2746 5704 2768
rect 1104 2694 1721 2746
rect 1773 2694 1785 2746
rect 1837 2694 1849 2746
rect 1901 2694 1913 2746
rect 1965 2694 1977 2746
rect 2029 2694 3262 2746
rect 3314 2694 3326 2746
rect 3378 2694 3390 2746
rect 3442 2694 3454 2746
rect 3506 2694 3518 2746
rect 3570 2694 4804 2746
rect 4856 2694 4868 2746
rect 4920 2694 4932 2746
rect 4984 2694 4996 2746
rect 5048 2694 5060 2746
rect 5112 2694 5704 2746
rect 1104 2672 5704 2694
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 2866 2428 2872 2440
rect 1719 2400 2872 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 4430 2388 4436 2440
rect 4488 2428 4494 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4488 2400 4721 2428
rect 4488 2388 4494 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1489 2295 1547 2301
rect 1489 2292 1501 2295
rect 72 2264 1501 2292
rect 72 2252 78 2264
rect 1489 2261 1501 2264
rect 1535 2261 1547 2295
rect 1489 2255 1547 2261
rect 4893 2295 4951 2301
rect 4893 2261 4905 2295
rect 4939 2292 4951 2295
rect 5810 2292 5816 2304
rect 4939 2264 5816 2292
rect 4939 2261 4951 2264
rect 4893 2255 4951 2261
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 1104 2202 5704 2224
rect 1104 2150 2491 2202
rect 2543 2150 2555 2202
rect 2607 2150 2619 2202
rect 2671 2150 2683 2202
rect 2735 2150 2747 2202
rect 2799 2150 4033 2202
rect 4085 2150 4097 2202
rect 4149 2150 4161 2202
rect 4213 2150 4225 2202
rect 4277 2150 4289 2202
rect 4341 2150 5704 2202
rect 1104 2128 5704 2150
<< via1 >>
rect 2491 8678 2543 8730
rect 2555 8678 2607 8730
rect 2619 8678 2671 8730
rect 2683 8678 2735 8730
rect 2747 8678 2799 8730
rect 4033 8678 4085 8730
rect 4097 8678 4149 8730
rect 4161 8678 4213 8730
rect 4225 8678 4277 8730
rect 4289 8678 4341 8730
rect 664 8576 716 8628
rect 6460 8576 6512 8628
rect 2136 8440 2188 8492
rect 4620 8440 4672 8492
rect 1721 8134 1773 8186
rect 1785 8134 1837 8186
rect 1849 8134 1901 8186
rect 1913 8134 1965 8186
rect 1977 8134 2029 8186
rect 3262 8134 3314 8186
rect 3326 8134 3378 8186
rect 3390 8134 3442 8186
rect 3454 8134 3506 8186
rect 3518 8134 3570 8186
rect 4804 8134 4856 8186
rect 4868 8134 4920 8186
rect 4932 8134 4984 8186
rect 4996 8134 5048 8186
rect 5060 8134 5112 8186
rect 2491 7590 2543 7642
rect 2555 7590 2607 7642
rect 2619 7590 2671 7642
rect 2683 7590 2735 7642
rect 2747 7590 2799 7642
rect 4033 7590 4085 7642
rect 4097 7590 4149 7642
rect 4161 7590 4213 7642
rect 4225 7590 4277 7642
rect 4289 7590 4341 7642
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 4436 7148 4488 7200
rect 1721 7046 1773 7098
rect 1785 7046 1837 7098
rect 1849 7046 1901 7098
rect 1913 7046 1965 7098
rect 1977 7046 2029 7098
rect 3262 7046 3314 7098
rect 3326 7046 3378 7098
rect 3390 7046 3442 7098
rect 3454 7046 3506 7098
rect 3518 7046 3570 7098
rect 4804 7046 4856 7098
rect 4868 7046 4920 7098
rect 4932 7046 4984 7098
rect 4996 7046 5048 7098
rect 5060 7046 5112 7098
rect 5172 6808 5224 6860
rect 2320 6740 2372 6792
rect 3884 6740 3936 6792
rect 4620 6740 4672 6792
rect 3700 6604 3752 6656
rect 4528 6604 4580 6656
rect 2491 6502 2543 6554
rect 2555 6502 2607 6554
rect 2619 6502 2671 6554
rect 2683 6502 2735 6554
rect 2747 6502 2799 6554
rect 4033 6502 4085 6554
rect 4097 6502 4149 6554
rect 4161 6502 4213 6554
rect 4225 6502 4277 6554
rect 4289 6502 4341 6554
rect 3608 6400 3660 6452
rect 3792 6332 3844 6384
rect 4620 6400 4672 6452
rect 1584 6264 1636 6316
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 4160 6239 4212 6248
rect 4160 6205 4169 6239
rect 4169 6205 4203 6239
rect 4203 6205 4212 6239
rect 4160 6196 4212 6205
rect 4528 6196 4580 6248
rect 2872 6060 2924 6112
rect 4528 6060 4580 6112
rect 1721 5958 1773 6010
rect 1785 5958 1837 6010
rect 1849 5958 1901 6010
rect 1913 5958 1965 6010
rect 1977 5958 2029 6010
rect 3262 5958 3314 6010
rect 3326 5958 3378 6010
rect 3390 5958 3442 6010
rect 3454 5958 3506 6010
rect 3518 5958 3570 6010
rect 4804 5958 4856 6010
rect 4868 5958 4920 6010
rect 4932 5958 4984 6010
rect 4996 5958 5048 6010
rect 5060 5958 5112 6010
rect 4160 5788 4212 5840
rect 3148 5652 3200 5704
rect 3700 5720 3752 5772
rect 4620 5720 4672 5772
rect 4436 5652 4488 5704
rect 5172 5652 5224 5704
rect 4712 5584 4764 5636
rect 2491 5414 2543 5466
rect 2555 5414 2607 5466
rect 2619 5414 2671 5466
rect 2683 5414 2735 5466
rect 2747 5414 2799 5466
rect 4033 5414 4085 5466
rect 4097 5414 4149 5466
rect 4161 5414 4213 5466
rect 4225 5414 4277 5466
rect 4289 5414 4341 5466
rect 2964 5287 3016 5296
rect 2964 5253 2973 5287
rect 2973 5253 3007 5287
rect 3007 5253 3016 5287
rect 2964 5244 3016 5253
rect 2228 5219 2280 5228
rect 2228 5185 2237 5219
rect 2237 5185 2271 5219
rect 2271 5185 2280 5219
rect 2228 5176 2280 5185
rect 3608 5108 3660 5160
rect 2136 4972 2188 5024
rect 3056 4972 3108 5024
rect 3884 4972 3936 5024
rect 1721 4870 1773 4922
rect 1785 4870 1837 4922
rect 1849 4870 1901 4922
rect 1913 4870 1965 4922
rect 1977 4870 2029 4922
rect 3262 4870 3314 4922
rect 3326 4870 3378 4922
rect 3390 4870 3442 4922
rect 3454 4870 3506 4922
rect 3518 4870 3570 4922
rect 4804 4870 4856 4922
rect 4868 4870 4920 4922
rect 4932 4870 4984 4922
rect 4996 4870 5048 4922
rect 5060 4870 5112 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 3056 4632 3108 4684
rect 4528 4700 4580 4752
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 3608 4564 3660 4616
rect 2044 4496 2096 4548
rect 3700 4496 3752 4548
rect 4436 4564 4488 4616
rect 5172 4564 5224 4616
rect 2491 4326 2543 4378
rect 2555 4326 2607 4378
rect 2619 4326 2671 4378
rect 2683 4326 2735 4378
rect 2747 4326 2799 4378
rect 4033 4326 4085 4378
rect 4097 4326 4149 4378
rect 4161 4326 4213 4378
rect 4225 4326 4277 4378
rect 4289 4326 4341 4378
rect 2044 4267 2096 4276
rect 2044 4233 2053 4267
rect 2053 4233 2087 4267
rect 2087 4233 2096 4267
rect 2044 4224 2096 4233
rect 2136 4088 2188 4140
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2872 4088 2924 4140
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 3700 4088 3752 4140
rect 4436 4088 4488 4140
rect 2964 4020 3016 4072
rect 3148 3952 3200 4004
rect 4528 3884 4580 3936
rect 1721 3782 1773 3834
rect 1785 3782 1837 3834
rect 1849 3782 1901 3834
rect 1913 3782 1965 3834
rect 1977 3782 2029 3834
rect 3262 3782 3314 3834
rect 3326 3782 3378 3834
rect 3390 3782 3442 3834
rect 3454 3782 3506 3834
rect 3518 3782 3570 3834
rect 4804 3782 4856 3834
rect 4868 3782 4920 3834
rect 4932 3782 4984 3834
rect 4996 3782 5048 3834
rect 5060 3782 5112 3834
rect 2964 3680 3016 3732
rect 3608 3680 3660 3732
rect 4436 3723 4488 3732
rect 4436 3689 4445 3723
rect 4445 3689 4479 3723
rect 4479 3689 4488 3723
rect 4436 3680 4488 3689
rect 2320 3544 2372 3596
rect 3884 3476 3936 3528
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4804 3476 4856 3528
rect 2491 3238 2543 3290
rect 2555 3238 2607 3290
rect 2619 3238 2671 3290
rect 2683 3238 2735 3290
rect 2747 3238 2799 3290
rect 4033 3238 4085 3290
rect 4097 3238 4149 3290
rect 4161 3238 4213 3290
rect 4225 3238 4277 3290
rect 4289 3238 4341 3290
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 5264 3000 5316 3052
rect 1721 2694 1773 2746
rect 1785 2694 1837 2746
rect 1849 2694 1901 2746
rect 1913 2694 1965 2746
rect 1977 2694 2029 2746
rect 3262 2694 3314 2746
rect 3326 2694 3378 2746
rect 3390 2694 3442 2746
rect 3454 2694 3506 2746
rect 3518 2694 3570 2746
rect 4804 2694 4856 2746
rect 4868 2694 4920 2746
rect 4932 2694 4984 2746
rect 4996 2694 5048 2746
rect 5060 2694 5112 2746
rect 2872 2388 2924 2440
rect 4436 2388 4488 2440
rect 20 2252 72 2304
rect 5816 2252 5868 2304
rect 2491 2150 2543 2202
rect 2555 2150 2607 2202
rect 2619 2150 2671 2202
rect 2683 2150 2735 2202
rect 2747 2150 2799 2202
rect 4033 2150 4085 2202
rect 4097 2150 4149 2202
rect 4161 2150 4213 2202
rect 4225 2150 4277 2202
rect 4289 2150 4341 2202
<< metal2 >>
rect 662 10177 718 10977
rect 6458 10177 6514 10977
rect 676 8634 704 10177
rect 2491 8732 2799 8752
rect 2491 8730 2497 8732
rect 2553 8730 2577 8732
rect 2633 8730 2657 8732
rect 2713 8730 2737 8732
rect 2793 8730 2799 8732
rect 2553 8678 2555 8730
rect 2735 8678 2737 8730
rect 2491 8676 2497 8678
rect 2553 8676 2577 8678
rect 2633 8676 2657 8678
rect 2713 8676 2737 8678
rect 2793 8676 2799 8678
rect 2491 8656 2799 8676
rect 4033 8732 4341 8752
rect 4033 8730 4039 8732
rect 4095 8730 4119 8732
rect 4175 8730 4199 8732
rect 4255 8730 4279 8732
rect 4335 8730 4341 8732
rect 4095 8678 4097 8730
rect 4277 8678 4279 8730
rect 4033 8676 4039 8678
rect 4095 8676 4119 8678
rect 4175 8676 4199 8678
rect 4255 8676 4279 8678
rect 4335 8676 4341 8678
rect 4033 8656 4341 8676
rect 6472 8634 6500 10177
rect 664 8628 716 8634
rect 664 8570 716 8576
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 1721 8188 2029 8208
rect 1721 8186 1727 8188
rect 1783 8186 1807 8188
rect 1863 8186 1887 8188
rect 1943 8186 1967 8188
rect 2023 8186 2029 8188
rect 1783 8134 1785 8186
rect 1965 8134 1967 8186
rect 1721 8132 1727 8134
rect 1783 8132 1807 8134
rect 1863 8132 1887 8134
rect 1943 8132 1967 8134
rect 2023 8132 2029 8134
rect 1721 8112 2029 8132
rect 1721 7100 2029 7120
rect 1721 7098 1727 7100
rect 1783 7098 1807 7100
rect 1863 7098 1887 7100
rect 1943 7098 1967 7100
rect 2023 7098 2029 7100
rect 1783 7046 1785 7098
rect 1965 7046 1967 7098
rect 1721 7044 1727 7046
rect 1783 7044 1807 7046
rect 1863 7044 1887 7046
rect 1943 7044 1967 7046
rect 2023 7044 2029 7046
rect 1721 7024 2029 7044
rect 2148 6322 2176 8434
rect 3262 8188 3570 8208
rect 3262 8186 3268 8188
rect 3324 8186 3348 8188
rect 3404 8186 3428 8188
rect 3484 8186 3508 8188
rect 3564 8186 3570 8188
rect 3324 8134 3326 8186
rect 3506 8134 3508 8186
rect 3262 8132 3268 8134
rect 3324 8132 3348 8134
rect 3404 8132 3428 8134
rect 3484 8132 3508 8134
rect 3564 8132 3570 8134
rect 3262 8112 3570 8132
rect 2491 7644 2799 7664
rect 2491 7642 2497 7644
rect 2553 7642 2577 7644
rect 2633 7642 2657 7644
rect 2713 7642 2737 7644
rect 2793 7642 2799 7644
rect 2553 7590 2555 7642
rect 2735 7590 2737 7642
rect 2491 7588 2497 7590
rect 2553 7588 2577 7590
rect 2633 7588 2657 7590
rect 2713 7588 2737 7590
rect 2793 7588 2799 7590
rect 2491 7568 2799 7588
rect 4033 7644 4341 7664
rect 4033 7642 4039 7644
rect 4095 7642 4119 7644
rect 4175 7642 4199 7644
rect 4255 7642 4279 7644
rect 4335 7642 4341 7644
rect 4095 7590 4097 7642
rect 4277 7590 4279 7642
rect 4033 7588 4039 7590
rect 4095 7588 4119 7590
rect 4175 7588 4199 7590
rect 4255 7588 4279 7590
rect 4335 7588 4341 7590
rect 4033 7568 4341 7588
rect 4632 7410 4660 8434
rect 4804 8188 5112 8208
rect 4804 8186 4810 8188
rect 4866 8186 4890 8188
rect 4946 8186 4970 8188
rect 5026 8186 5050 8188
rect 5106 8186 5112 8188
rect 4866 8134 4868 8186
rect 5048 8134 5050 8186
rect 4804 8132 4810 8134
rect 4866 8132 4890 8134
rect 4946 8132 4970 8134
rect 5026 8132 5050 8134
rect 5106 8132 5112 8134
rect 4804 8112 5112 8132
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 3262 7100 3570 7120
rect 3262 7098 3268 7100
rect 3324 7098 3348 7100
rect 3404 7098 3428 7100
rect 3484 7098 3508 7100
rect 3564 7098 3570 7100
rect 3324 7046 3326 7098
rect 3506 7046 3508 7098
rect 3262 7044 3268 7046
rect 3324 7044 3348 7046
rect 3404 7044 3428 7046
rect 3484 7044 3508 7046
rect 3564 7044 3570 7046
rect 3262 7024 3570 7044
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 1596 4826 1624 6258
rect 1721 6012 2029 6032
rect 1721 6010 1727 6012
rect 1783 6010 1807 6012
rect 1863 6010 1887 6012
rect 1943 6010 1967 6012
rect 2023 6010 2029 6012
rect 1783 5958 1785 6010
rect 1965 5958 1967 6010
rect 1721 5956 1727 5958
rect 1783 5956 1807 5958
rect 1863 5956 1887 5958
rect 1943 5956 1967 5958
rect 2023 5956 2029 5958
rect 1721 5936 2029 5956
rect 2240 5234 2268 6258
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 1721 4924 2029 4944
rect 1721 4922 1727 4924
rect 1783 4922 1807 4924
rect 1863 4922 1887 4924
rect 1943 4922 1967 4924
rect 2023 4922 2029 4924
rect 1783 4870 1785 4922
rect 1965 4870 1967 4922
rect 1721 4868 1727 4870
rect 1783 4868 1807 4870
rect 1863 4868 1887 4870
rect 1943 4868 1967 4870
rect 2023 4868 2029 4870
rect 1721 4848 2029 4868
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 2044 4548 2096 4554
rect 2044 4490 2096 4496
rect 2056 4282 2084 4490
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 2148 4146 2176 4966
rect 2332 4146 2360 6734
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 2491 6556 2799 6576
rect 2491 6554 2497 6556
rect 2553 6554 2577 6556
rect 2633 6554 2657 6556
rect 2713 6554 2737 6556
rect 2793 6554 2799 6556
rect 2553 6502 2555 6554
rect 2735 6502 2737 6554
rect 2491 6500 2497 6502
rect 2553 6500 2577 6502
rect 2633 6500 2657 6502
rect 2713 6500 2737 6502
rect 2793 6500 2799 6502
rect 2491 6480 2799 6500
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2491 5468 2799 5488
rect 2491 5466 2497 5468
rect 2553 5466 2577 5468
rect 2633 5466 2657 5468
rect 2713 5466 2737 5468
rect 2793 5466 2799 5468
rect 2553 5414 2555 5466
rect 2735 5414 2737 5466
rect 2491 5412 2497 5414
rect 2553 5412 2577 5414
rect 2633 5412 2657 5414
rect 2713 5412 2737 5414
rect 2793 5412 2799 5414
rect 2491 5392 2799 5412
rect 2491 4380 2799 4400
rect 2491 4378 2497 4380
rect 2553 4378 2577 4380
rect 2633 4378 2657 4380
rect 2713 4378 2737 4380
rect 2793 4378 2799 4380
rect 2553 4326 2555 4378
rect 2735 4326 2737 4378
rect 2491 4324 2497 4326
rect 2553 4324 2577 4326
rect 2633 4324 2657 4326
rect 2713 4324 2737 4326
rect 2793 4324 2799 4326
rect 2491 4304 2799 4324
rect 2884 4146 2912 6054
rect 3262 6012 3570 6032
rect 3262 6010 3268 6012
rect 3324 6010 3348 6012
rect 3404 6010 3428 6012
rect 3484 6010 3508 6012
rect 3564 6010 3570 6012
rect 3324 5958 3326 6010
rect 3506 5958 3508 6010
rect 3262 5956 3268 5958
rect 3324 5956 3348 5958
rect 3404 5956 3428 5958
rect 3484 5956 3508 5958
rect 3564 5956 3570 5958
rect 3262 5936 3570 5956
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2964 5296 3016 5302
rect 2962 5264 2964 5273
rect 3016 5264 3018 5273
rect 2962 5199 3018 5208
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3068 4690 3096 4966
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 1721 3836 2029 3856
rect 1721 3834 1727 3836
rect 1783 3834 1807 3836
rect 1863 3834 1887 3836
rect 1943 3834 1967 3836
rect 2023 3834 2029 3836
rect 1783 3782 1785 3834
rect 1965 3782 1967 3834
rect 1721 3780 1727 3782
rect 1783 3780 1807 3782
rect 1863 3780 1887 3782
rect 1943 3780 1967 3782
rect 2023 3780 2029 3782
rect 1721 3760 2029 3780
rect 2332 3602 2360 4082
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2491 3292 2799 3312
rect 2491 3290 2497 3292
rect 2553 3290 2577 3292
rect 2633 3290 2657 3292
rect 2713 3290 2737 3292
rect 2793 3290 2799 3292
rect 2553 3238 2555 3290
rect 2735 3238 2737 3290
rect 2491 3236 2497 3238
rect 2553 3236 2577 3238
rect 2633 3236 2657 3238
rect 2713 3236 2737 3238
rect 2793 3236 2799 3238
rect 2491 3216 2799 3236
rect 1721 2748 2029 2768
rect 1721 2746 1727 2748
rect 1783 2746 1807 2748
rect 1863 2746 1887 2748
rect 1943 2746 1967 2748
rect 2023 2746 2029 2748
rect 1783 2694 1785 2746
rect 1965 2694 1967 2746
rect 1721 2692 1727 2694
rect 1783 2692 1807 2694
rect 1863 2692 1887 2694
rect 1943 2692 1967 2694
rect 2023 2692 2029 2694
rect 1721 2672 2029 2692
rect 2884 2446 2912 4082
rect 2976 4078 3004 4558
rect 3068 4146 3096 4626
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2976 3738 3004 4014
rect 3160 4010 3188 5646
rect 3620 5166 3648 6394
rect 3712 5778 3740 6598
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3262 4924 3570 4944
rect 3262 4922 3268 4924
rect 3324 4922 3348 4924
rect 3404 4922 3428 4924
rect 3484 4922 3508 4924
rect 3564 4922 3570 4924
rect 3324 4870 3326 4922
rect 3506 4870 3508 4922
rect 3262 4868 3268 4870
rect 3324 4868 3348 4870
rect 3404 4868 3428 4870
rect 3484 4868 3508 4870
rect 3564 4868 3570 4870
rect 3262 4848 3570 4868
rect 3620 4622 3648 5102
rect 3804 4826 3832 6326
rect 3896 5030 3924 6734
rect 4033 6556 4341 6576
rect 4033 6554 4039 6556
rect 4095 6554 4119 6556
rect 4175 6554 4199 6556
rect 4255 6554 4279 6556
rect 4335 6554 4341 6556
rect 4095 6502 4097 6554
rect 4277 6502 4279 6554
rect 4033 6500 4039 6502
rect 4095 6500 4119 6502
rect 4175 6500 4199 6502
rect 4255 6500 4279 6502
rect 4335 6500 4341 6502
rect 4033 6480 4341 6500
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4172 5846 4200 6190
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 4448 5710 4476 7142
rect 4632 6914 4660 7346
rect 4804 7100 5112 7120
rect 4804 7098 4810 7100
rect 4866 7098 4890 7100
rect 4946 7098 4970 7100
rect 5026 7098 5050 7100
rect 5106 7098 5112 7100
rect 4866 7046 4868 7098
rect 5048 7046 5050 7098
rect 4804 7044 4810 7046
rect 4866 7044 4890 7046
rect 4946 7044 4970 7046
rect 5026 7044 5050 7046
rect 5106 7044 5112 7046
rect 4804 7024 5112 7044
rect 4632 6886 4752 6914
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6254 4568 6598
rect 4632 6458 4660 6734
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4033 5468 4341 5488
rect 4033 5466 4039 5468
rect 4095 5466 4119 5468
rect 4175 5466 4199 5468
rect 4255 5466 4279 5468
rect 4335 5466 4341 5468
rect 4095 5414 4097 5466
rect 4277 5414 4279 5466
rect 4033 5412 4039 5414
rect 4095 5412 4119 5414
rect 4175 5412 4199 5414
rect 4255 5412 4279 5414
rect 4335 5412 4341 5414
rect 4033 5392 4341 5412
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3262 3836 3570 3856
rect 3262 3834 3268 3836
rect 3324 3834 3348 3836
rect 3404 3834 3428 3836
rect 3484 3834 3508 3836
rect 3564 3834 3570 3836
rect 3324 3782 3326 3834
rect 3506 3782 3508 3834
rect 3262 3780 3268 3782
rect 3324 3780 3348 3782
rect 3404 3780 3428 3782
rect 3484 3780 3508 3782
rect 3564 3780 3570 3782
rect 3262 3760 3570 3780
rect 3620 3738 3648 4558
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3712 4146 3740 4490
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3896 3534 3924 4966
rect 4540 4758 4568 6054
rect 4632 5778 4660 6394
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4724 5642 4752 6886
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 4804 6012 5112 6032
rect 4804 6010 4810 6012
rect 4866 6010 4890 6012
rect 4946 6010 4970 6012
rect 5026 6010 5050 6012
rect 5106 6010 5112 6012
rect 4866 5958 4868 6010
rect 5048 5958 5050 6010
rect 4804 5956 4810 5958
rect 4866 5956 4890 5958
rect 4946 5956 4970 5958
rect 5026 5956 5050 5958
rect 5106 5956 5112 5958
rect 4804 5936 5112 5956
rect 5184 5710 5212 6802
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4804 4924 5112 4944
rect 4804 4922 4810 4924
rect 4866 4922 4890 4924
rect 4946 4922 4970 4924
rect 5026 4922 5050 4924
rect 5106 4922 5112 4924
rect 4866 4870 4868 4922
rect 5048 4870 5050 4922
rect 4804 4868 4810 4870
rect 4866 4868 4890 4870
rect 4946 4868 4970 4870
rect 5026 4868 5050 4870
rect 5106 4868 5112 4870
rect 4804 4848 5112 4868
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 5184 4622 5212 5646
rect 5262 4856 5318 4865
rect 5262 4791 5318 4800
rect 4436 4616 4488 4622
rect 5172 4616 5224 4622
rect 4488 4564 4568 4570
rect 4436 4558 4568 4564
rect 5172 4558 5224 4564
rect 4448 4542 4568 4558
rect 4033 4380 4341 4400
rect 4033 4378 4039 4380
rect 4095 4378 4119 4380
rect 4175 4378 4199 4380
rect 4255 4378 4279 4380
rect 4335 4378 4341 4380
rect 4095 4326 4097 4378
rect 4277 4326 4279 4378
rect 4033 4324 4039 4326
rect 4095 4324 4119 4326
rect 4175 4324 4199 4326
rect 4255 4324 4279 4326
rect 4335 4324 4341 4326
rect 4033 4304 4341 4324
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4448 3738 4476 4082
rect 4540 3942 4568 4542
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4540 3618 4568 3878
rect 4804 3836 5112 3856
rect 4804 3834 4810 3836
rect 4866 3834 4890 3836
rect 4946 3834 4970 3836
rect 5026 3834 5050 3836
rect 5106 3834 5112 3836
rect 4866 3782 4868 3834
rect 5048 3782 5050 3834
rect 4804 3780 4810 3782
rect 4866 3780 4890 3782
rect 4946 3780 4970 3782
rect 5026 3780 5050 3782
rect 5106 3780 5112 3782
rect 4804 3760 5112 3780
rect 4448 3590 4568 3618
rect 4448 3534 4476 3590
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4033 3292 4341 3312
rect 4033 3290 4039 3292
rect 4095 3290 4119 3292
rect 4175 3290 4199 3292
rect 4255 3290 4279 3292
rect 4335 3290 4341 3292
rect 4095 3238 4097 3290
rect 4277 3238 4279 3290
rect 4033 3236 4039 3238
rect 4095 3236 4119 3238
rect 4175 3236 4199 3238
rect 4255 3236 4279 3238
rect 4335 3236 4341 3238
rect 4033 3216 4341 3236
rect 3262 2748 3570 2768
rect 3262 2746 3268 2748
rect 3324 2746 3348 2748
rect 3404 2746 3428 2748
rect 3484 2746 3508 2748
rect 3564 2746 3570 2748
rect 3324 2694 3326 2746
rect 3506 2694 3508 2746
rect 3262 2692 3268 2694
rect 3324 2692 3348 2694
rect 3404 2692 3428 2694
rect 3484 2692 3508 2694
rect 3564 2692 3570 2694
rect 3262 2672 3570 2692
rect 4448 2446 4476 3470
rect 4816 3194 4844 3470
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5276 3058 5304 4791
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 4804 2748 5112 2768
rect 4804 2746 4810 2748
rect 4866 2746 4890 2748
rect 4946 2746 4970 2748
rect 5026 2746 5050 2748
rect 5106 2746 5112 2748
rect 4866 2694 4868 2746
rect 5048 2694 5050 2746
rect 4804 2692 4810 2694
rect 4866 2692 4890 2694
rect 4946 2692 4970 2694
rect 5026 2692 5050 2694
rect 5106 2692 5112 2694
rect 4804 2672 5112 2692
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 32 800 60 2246
rect 2491 2204 2799 2224
rect 2491 2202 2497 2204
rect 2553 2202 2577 2204
rect 2633 2202 2657 2204
rect 2713 2202 2737 2204
rect 2793 2202 2799 2204
rect 2553 2150 2555 2202
rect 2735 2150 2737 2202
rect 2491 2148 2497 2150
rect 2553 2148 2577 2150
rect 2633 2148 2657 2150
rect 2713 2148 2737 2150
rect 2793 2148 2799 2150
rect 2491 2128 2799 2148
rect 4033 2204 4341 2224
rect 4033 2202 4039 2204
rect 4095 2202 4119 2204
rect 4175 2202 4199 2204
rect 4255 2202 4279 2204
rect 4335 2202 4341 2204
rect 4095 2150 4097 2202
rect 4277 2150 4279 2202
rect 4033 2148 4039 2150
rect 4095 2148 4119 2150
rect 4175 2148 4199 2150
rect 4255 2148 4279 2150
rect 4335 2148 4341 2150
rect 4033 2128 4341 2148
rect 5828 800 5856 2246
rect 18 0 74 800
rect 5814 0 5870 800
<< via2 >>
rect 2497 8730 2553 8732
rect 2577 8730 2633 8732
rect 2657 8730 2713 8732
rect 2737 8730 2793 8732
rect 2497 8678 2543 8730
rect 2543 8678 2553 8730
rect 2577 8678 2607 8730
rect 2607 8678 2619 8730
rect 2619 8678 2633 8730
rect 2657 8678 2671 8730
rect 2671 8678 2683 8730
rect 2683 8678 2713 8730
rect 2737 8678 2747 8730
rect 2747 8678 2793 8730
rect 2497 8676 2553 8678
rect 2577 8676 2633 8678
rect 2657 8676 2713 8678
rect 2737 8676 2793 8678
rect 4039 8730 4095 8732
rect 4119 8730 4175 8732
rect 4199 8730 4255 8732
rect 4279 8730 4335 8732
rect 4039 8678 4085 8730
rect 4085 8678 4095 8730
rect 4119 8678 4149 8730
rect 4149 8678 4161 8730
rect 4161 8678 4175 8730
rect 4199 8678 4213 8730
rect 4213 8678 4225 8730
rect 4225 8678 4255 8730
rect 4279 8678 4289 8730
rect 4289 8678 4335 8730
rect 4039 8676 4095 8678
rect 4119 8676 4175 8678
rect 4199 8676 4255 8678
rect 4279 8676 4335 8678
rect 1727 8186 1783 8188
rect 1807 8186 1863 8188
rect 1887 8186 1943 8188
rect 1967 8186 2023 8188
rect 1727 8134 1773 8186
rect 1773 8134 1783 8186
rect 1807 8134 1837 8186
rect 1837 8134 1849 8186
rect 1849 8134 1863 8186
rect 1887 8134 1901 8186
rect 1901 8134 1913 8186
rect 1913 8134 1943 8186
rect 1967 8134 1977 8186
rect 1977 8134 2023 8186
rect 1727 8132 1783 8134
rect 1807 8132 1863 8134
rect 1887 8132 1943 8134
rect 1967 8132 2023 8134
rect 1727 7098 1783 7100
rect 1807 7098 1863 7100
rect 1887 7098 1943 7100
rect 1967 7098 2023 7100
rect 1727 7046 1773 7098
rect 1773 7046 1783 7098
rect 1807 7046 1837 7098
rect 1837 7046 1849 7098
rect 1849 7046 1863 7098
rect 1887 7046 1901 7098
rect 1901 7046 1913 7098
rect 1913 7046 1943 7098
rect 1967 7046 1977 7098
rect 1977 7046 2023 7098
rect 1727 7044 1783 7046
rect 1807 7044 1863 7046
rect 1887 7044 1943 7046
rect 1967 7044 2023 7046
rect 3268 8186 3324 8188
rect 3348 8186 3404 8188
rect 3428 8186 3484 8188
rect 3508 8186 3564 8188
rect 3268 8134 3314 8186
rect 3314 8134 3324 8186
rect 3348 8134 3378 8186
rect 3378 8134 3390 8186
rect 3390 8134 3404 8186
rect 3428 8134 3442 8186
rect 3442 8134 3454 8186
rect 3454 8134 3484 8186
rect 3508 8134 3518 8186
rect 3518 8134 3564 8186
rect 3268 8132 3324 8134
rect 3348 8132 3404 8134
rect 3428 8132 3484 8134
rect 3508 8132 3564 8134
rect 2497 7642 2553 7644
rect 2577 7642 2633 7644
rect 2657 7642 2713 7644
rect 2737 7642 2793 7644
rect 2497 7590 2543 7642
rect 2543 7590 2553 7642
rect 2577 7590 2607 7642
rect 2607 7590 2619 7642
rect 2619 7590 2633 7642
rect 2657 7590 2671 7642
rect 2671 7590 2683 7642
rect 2683 7590 2713 7642
rect 2737 7590 2747 7642
rect 2747 7590 2793 7642
rect 2497 7588 2553 7590
rect 2577 7588 2633 7590
rect 2657 7588 2713 7590
rect 2737 7588 2793 7590
rect 4039 7642 4095 7644
rect 4119 7642 4175 7644
rect 4199 7642 4255 7644
rect 4279 7642 4335 7644
rect 4039 7590 4085 7642
rect 4085 7590 4095 7642
rect 4119 7590 4149 7642
rect 4149 7590 4161 7642
rect 4161 7590 4175 7642
rect 4199 7590 4213 7642
rect 4213 7590 4225 7642
rect 4225 7590 4255 7642
rect 4279 7590 4289 7642
rect 4289 7590 4335 7642
rect 4039 7588 4095 7590
rect 4119 7588 4175 7590
rect 4199 7588 4255 7590
rect 4279 7588 4335 7590
rect 4810 8186 4866 8188
rect 4890 8186 4946 8188
rect 4970 8186 5026 8188
rect 5050 8186 5106 8188
rect 4810 8134 4856 8186
rect 4856 8134 4866 8186
rect 4890 8134 4920 8186
rect 4920 8134 4932 8186
rect 4932 8134 4946 8186
rect 4970 8134 4984 8186
rect 4984 8134 4996 8186
rect 4996 8134 5026 8186
rect 5050 8134 5060 8186
rect 5060 8134 5106 8186
rect 4810 8132 4866 8134
rect 4890 8132 4946 8134
rect 4970 8132 5026 8134
rect 5050 8132 5106 8134
rect 3268 7098 3324 7100
rect 3348 7098 3404 7100
rect 3428 7098 3484 7100
rect 3508 7098 3564 7100
rect 3268 7046 3314 7098
rect 3314 7046 3324 7098
rect 3348 7046 3378 7098
rect 3378 7046 3390 7098
rect 3390 7046 3404 7098
rect 3428 7046 3442 7098
rect 3442 7046 3454 7098
rect 3454 7046 3484 7098
rect 3508 7046 3518 7098
rect 3518 7046 3564 7098
rect 3268 7044 3324 7046
rect 3348 7044 3404 7046
rect 3428 7044 3484 7046
rect 3508 7044 3564 7046
rect 1727 6010 1783 6012
rect 1807 6010 1863 6012
rect 1887 6010 1943 6012
rect 1967 6010 2023 6012
rect 1727 5958 1773 6010
rect 1773 5958 1783 6010
rect 1807 5958 1837 6010
rect 1837 5958 1849 6010
rect 1849 5958 1863 6010
rect 1887 5958 1901 6010
rect 1901 5958 1913 6010
rect 1913 5958 1943 6010
rect 1967 5958 1977 6010
rect 1977 5958 2023 6010
rect 1727 5956 1783 5958
rect 1807 5956 1863 5958
rect 1887 5956 1943 5958
rect 1967 5956 2023 5958
rect 1727 4922 1783 4924
rect 1807 4922 1863 4924
rect 1887 4922 1943 4924
rect 1967 4922 2023 4924
rect 1727 4870 1773 4922
rect 1773 4870 1783 4922
rect 1807 4870 1837 4922
rect 1837 4870 1849 4922
rect 1849 4870 1863 4922
rect 1887 4870 1901 4922
rect 1901 4870 1913 4922
rect 1913 4870 1943 4922
rect 1967 4870 1977 4922
rect 1977 4870 2023 4922
rect 1727 4868 1783 4870
rect 1807 4868 1863 4870
rect 1887 4868 1943 4870
rect 1967 4868 2023 4870
rect 2497 6554 2553 6556
rect 2577 6554 2633 6556
rect 2657 6554 2713 6556
rect 2737 6554 2793 6556
rect 2497 6502 2543 6554
rect 2543 6502 2553 6554
rect 2577 6502 2607 6554
rect 2607 6502 2619 6554
rect 2619 6502 2633 6554
rect 2657 6502 2671 6554
rect 2671 6502 2683 6554
rect 2683 6502 2713 6554
rect 2737 6502 2747 6554
rect 2747 6502 2793 6554
rect 2497 6500 2553 6502
rect 2577 6500 2633 6502
rect 2657 6500 2713 6502
rect 2737 6500 2793 6502
rect 2497 5466 2553 5468
rect 2577 5466 2633 5468
rect 2657 5466 2713 5468
rect 2737 5466 2793 5468
rect 2497 5414 2543 5466
rect 2543 5414 2553 5466
rect 2577 5414 2607 5466
rect 2607 5414 2619 5466
rect 2619 5414 2633 5466
rect 2657 5414 2671 5466
rect 2671 5414 2683 5466
rect 2683 5414 2713 5466
rect 2737 5414 2747 5466
rect 2747 5414 2793 5466
rect 2497 5412 2553 5414
rect 2577 5412 2633 5414
rect 2657 5412 2713 5414
rect 2737 5412 2793 5414
rect 2497 4378 2553 4380
rect 2577 4378 2633 4380
rect 2657 4378 2713 4380
rect 2737 4378 2793 4380
rect 2497 4326 2543 4378
rect 2543 4326 2553 4378
rect 2577 4326 2607 4378
rect 2607 4326 2619 4378
rect 2619 4326 2633 4378
rect 2657 4326 2671 4378
rect 2671 4326 2683 4378
rect 2683 4326 2713 4378
rect 2737 4326 2747 4378
rect 2747 4326 2793 4378
rect 2497 4324 2553 4326
rect 2577 4324 2633 4326
rect 2657 4324 2713 4326
rect 2737 4324 2793 4326
rect 3268 6010 3324 6012
rect 3348 6010 3404 6012
rect 3428 6010 3484 6012
rect 3508 6010 3564 6012
rect 3268 5958 3314 6010
rect 3314 5958 3324 6010
rect 3348 5958 3378 6010
rect 3378 5958 3390 6010
rect 3390 5958 3404 6010
rect 3428 5958 3442 6010
rect 3442 5958 3454 6010
rect 3454 5958 3484 6010
rect 3508 5958 3518 6010
rect 3518 5958 3564 6010
rect 3268 5956 3324 5958
rect 3348 5956 3404 5958
rect 3428 5956 3484 5958
rect 3508 5956 3564 5958
rect 2962 5244 2964 5264
rect 2964 5244 3016 5264
rect 3016 5244 3018 5264
rect 2962 5208 3018 5244
rect 1727 3834 1783 3836
rect 1807 3834 1863 3836
rect 1887 3834 1943 3836
rect 1967 3834 2023 3836
rect 1727 3782 1773 3834
rect 1773 3782 1783 3834
rect 1807 3782 1837 3834
rect 1837 3782 1849 3834
rect 1849 3782 1863 3834
rect 1887 3782 1901 3834
rect 1901 3782 1913 3834
rect 1913 3782 1943 3834
rect 1967 3782 1977 3834
rect 1977 3782 2023 3834
rect 1727 3780 1783 3782
rect 1807 3780 1863 3782
rect 1887 3780 1943 3782
rect 1967 3780 2023 3782
rect 2497 3290 2553 3292
rect 2577 3290 2633 3292
rect 2657 3290 2713 3292
rect 2737 3290 2793 3292
rect 2497 3238 2543 3290
rect 2543 3238 2553 3290
rect 2577 3238 2607 3290
rect 2607 3238 2619 3290
rect 2619 3238 2633 3290
rect 2657 3238 2671 3290
rect 2671 3238 2683 3290
rect 2683 3238 2713 3290
rect 2737 3238 2747 3290
rect 2747 3238 2793 3290
rect 2497 3236 2553 3238
rect 2577 3236 2633 3238
rect 2657 3236 2713 3238
rect 2737 3236 2793 3238
rect 1727 2746 1783 2748
rect 1807 2746 1863 2748
rect 1887 2746 1943 2748
rect 1967 2746 2023 2748
rect 1727 2694 1773 2746
rect 1773 2694 1783 2746
rect 1807 2694 1837 2746
rect 1837 2694 1849 2746
rect 1849 2694 1863 2746
rect 1887 2694 1901 2746
rect 1901 2694 1913 2746
rect 1913 2694 1943 2746
rect 1967 2694 1977 2746
rect 1977 2694 2023 2746
rect 1727 2692 1783 2694
rect 1807 2692 1863 2694
rect 1887 2692 1943 2694
rect 1967 2692 2023 2694
rect 3268 4922 3324 4924
rect 3348 4922 3404 4924
rect 3428 4922 3484 4924
rect 3508 4922 3564 4924
rect 3268 4870 3314 4922
rect 3314 4870 3324 4922
rect 3348 4870 3378 4922
rect 3378 4870 3390 4922
rect 3390 4870 3404 4922
rect 3428 4870 3442 4922
rect 3442 4870 3454 4922
rect 3454 4870 3484 4922
rect 3508 4870 3518 4922
rect 3518 4870 3564 4922
rect 3268 4868 3324 4870
rect 3348 4868 3404 4870
rect 3428 4868 3484 4870
rect 3508 4868 3564 4870
rect 4039 6554 4095 6556
rect 4119 6554 4175 6556
rect 4199 6554 4255 6556
rect 4279 6554 4335 6556
rect 4039 6502 4085 6554
rect 4085 6502 4095 6554
rect 4119 6502 4149 6554
rect 4149 6502 4161 6554
rect 4161 6502 4175 6554
rect 4199 6502 4213 6554
rect 4213 6502 4225 6554
rect 4225 6502 4255 6554
rect 4279 6502 4289 6554
rect 4289 6502 4335 6554
rect 4039 6500 4095 6502
rect 4119 6500 4175 6502
rect 4199 6500 4255 6502
rect 4279 6500 4335 6502
rect 4810 7098 4866 7100
rect 4890 7098 4946 7100
rect 4970 7098 5026 7100
rect 5050 7098 5106 7100
rect 4810 7046 4856 7098
rect 4856 7046 4866 7098
rect 4890 7046 4920 7098
rect 4920 7046 4932 7098
rect 4932 7046 4946 7098
rect 4970 7046 4984 7098
rect 4984 7046 4996 7098
rect 4996 7046 5026 7098
rect 5050 7046 5060 7098
rect 5060 7046 5106 7098
rect 4810 7044 4866 7046
rect 4890 7044 4946 7046
rect 4970 7044 5026 7046
rect 5050 7044 5106 7046
rect 4039 5466 4095 5468
rect 4119 5466 4175 5468
rect 4199 5466 4255 5468
rect 4279 5466 4335 5468
rect 4039 5414 4085 5466
rect 4085 5414 4095 5466
rect 4119 5414 4149 5466
rect 4149 5414 4161 5466
rect 4161 5414 4175 5466
rect 4199 5414 4213 5466
rect 4213 5414 4225 5466
rect 4225 5414 4255 5466
rect 4279 5414 4289 5466
rect 4289 5414 4335 5466
rect 4039 5412 4095 5414
rect 4119 5412 4175 5414
rect 4199 5412 4255 5414
rect 4279 5412 4335 5414
rect 3268 3834 3324 3836
rect 3348 3834 3404 3836
rect 3428 3834 3484 3836
rect 3508 3834 3564 3836
rect 3268 3782 3314 3834
rect 3314 3782 3324 3834
rect 3348 3782 3378 3834
rect 3378 3782 3390 3834
rect 3390 3782 3404 3834
rect 3428 3782 3442 3834
rect 3442 3782 3454 3834
rect 3454 3782 3484 3834
rect 3508 3782 3518 3834
rect 3518 3782 3564 3834
rect 3268 3780 3324 3782
rect 3348 3780 3404 3782
rect 3428 3780 3484 3782
rect 3508 3780 3564 3782
rect 4810 6010 4866 6012
rect 4890 6010 4946 6012
rect 4970 6010 5026 6012
rect 5050 6010 5106 6012
rect 4810 5958 4856 6010
rect 4856 5958 4866 6010
rect 4890 5958 4920 6010
rect 4920 5958 4932 6010
rect 4932 5958 4946 6010
rect 4970 5958 4984 6010
rect 4984 5958 4996 6010
rect 4996 5958 5026 6010
rect 5050 5958 5060 6010
rect 5060 5958 5106 6010
rect 4810 5956 4866 5958
rect 4890 5956 4946 5958
rect 4970 5956 5026 5958
rect 5050 5956 5106 5958
rect 4810 4922 4866 4924
rect 4890 4922 4946 4924
rect 4970 4922 5026 4924
rect 5050 4922 5106 4924
rect 4810 4870 4856 4922
rect 4856 4870 4866 4922
rect 4890 4870 4920 4922
rect 4920 4870 4932 4922
rect 4932 4870 4946 4922
rect 4970 4870 4984 4922
rect 4984 4870 4996 4922
rect 4996 4870 5026 4922
rect 5050 4870 5060 4922
rect 5060 4870 5106 4922
rect 4810 4868 4866 4870
rect 4890 4868 4946 4870
rect 4970 4868 5026 4870
rect 5050 4868 5106 4870
rect 5262 4800 5318 4856
rect 4039 4378 4095 4380
rect 4119 4378 4175 4380
rect 4199 4378 4255 4380
rect 4279 4378 4335 4380
rect 4039 4326 4085 4378
rect 4085 4326 4095 4378
rect 4119 4326 4149 4378
rect 4149 4326 4161 4378
rect 4161 4326 4175 4378
rect 4199 4326 4213 4378
rect 4213 4326 4225 4378
rect 4225 4326 4255 4378
rect 4279 4326 4289 4378
rect 4289 4326 4335 4378
rect 4039 4324 4095 4326
rect 4119 4324 4175 4326
rect 4199 4324 4255 4326
rect 4279 4324 4335 4326
rect 4810 3834 4866 3836
rect 4890 3834 4946 3836
rect 4970 3834 5026 3836
rect 5050 3834 5106 3836
rect 4810 3782 4856 3834
rect 4856 3782 4866 3834
rect 4890 3782 4920 3834
rect 4920 3782 4932 3834
rect 4932 3782 4946 3834
rect 4970 3782 4984 3834
rect 4984 3782 4996 3834
rect 4996 3782 5026 3834
rect 5050 3782 5060 3834
rect 5060 3782 5106 3834
rect 4810 3780 4866 3782
rect 4890 3780 4946 3782
rect 4970 3780 5026 3782
rect 5050 3780 5106 3782
rect 4039 3290 4095 3292
rect 4119 3290 4175 3292
rect 4199 3290 4255 3292
rect 4279 3290 4335 3292
rect 4039 3238 4085 3290
rect 4085 3238 4095 3290
rect 4119 3238 4149 3290
rect 4149 3238 4161 3290
rect 4161 3238 4175 3290
rect 4199 3238 4213 3290
rect 4213 3238 4225 3290
rect 4225 3238 4255 3290
rect 4279 3238 4289 3290
rect 4289 3238 4335 3290
rect 4039 3236 4095 3238
rect 4119 3236 4175 3238
rect 4199 3236 4255 3238
rect 4279 3236 4335 3238
rect 3268 2746 3324 2748
rect 3348 2746 3404 2748
rect 3428 2746 3484 2748
rect 3508 2746 3564 2748
rect 3268 2694 3314 2746
rect 3314 2694 3324 2746
rect 3348 2694 3378 2746
rect 3378 2694 3390 2746
rect 3390 2694 3404 2746
rect 3428 2694 3442 2746
rect 3442 2694 3454 2746
rect 3454 2694 3484 2746
rect 3508 2694 3518 2746
rect 3518 2694 3564 2746
rect 3268 2692 3324 2694
rect 3348 2692 3404 2694
rect 3428 2692 3484 2694
rect 3508 2692 3564 2694
rect 4810 2746 4866 2748
rect 4890 2746 4946 2748
rect 4970 2746 5026 2748
rect 5050 2746 5106 2748
rect 4810 2694 4856 2746
rect 4856 2694 4866 2746
rect 4890 2694 4920 2746
rect 4920 2694 4932 2746
rect 4932 2694 4946 2746
rect 4970 2694 4984 2746
rect 4984 2694 4996 2746
rect 4996 2694 5026 2746
rect 5050 2694 5060 2746
rect 5060 2694 5106 2746
rect 4810 2692 4866 2694
rect 4890 2692 4946 2694
rect 4970 2692 5026 2694
rect 5050 2692 5106 2694
rect 2497 2202 2553 2204
rect 2577 2202 2633 2204
rect 2657 2202 2713 2204
rect 2737 2202 2793 2204
rect 2497 2150 2543 2202
rect 2543 2150 2553 2202
rect 2577 2150 2607 2202
rect 2607 2150 2619 2202
rect 2619 2150 2633 2202
rect 2657 2150 2671 2202
rect 2671 2150 2683 2202
rect 2683 2150 2713 2202
rect 2737 2150 2747 2202
rect 2747 2150 2793 2202
rect 2497 2148 2553 2150
rect 2577 2148 2633 2150
rect 2657 2148 2713 2150
rect 2737 2148 2793 2150
rect 4039 2202 4095 2204
rect 4119 2202 4175 2204
rect 4199 2202 4255 2204
rect 4279 2202 4335 2204
rect 4039 2150 4085 2202
rect 4085 2150 4095 2202
rect 4119 2150 4149 2202
rect 4149 2150 4161 2202
rect 4161 2150 4175 2202
rect 4199 2150 4213 2202
rect 4213 2150 4225 2202
rect 4225 2150 4255 2202
rect 4279 2150 4289 2202
rect 4289 2150 4335 2202
rect 4039 2148 4095 2150
rect 4119 2148 4175 2150
rect 4199 2148 4255 2150
rect 4279 2148 4335 2150
<< metal3 >>
rect 2485 8736 2805 8737
rect 2485 8672 2493 8736
rect 2557 8672 2573 8736
rect 2637 8672 2653 8736
rect 2717 8672 2733 8736
rect 2797 8672 2805 8736
rect 2485 8671 2805 8672
rect 4027 8736 4347 8737
rect 4027 8672 4035 8736
rect 4099 8672 4115 8736
rect 4179 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4347 8736
rect 4027 8671 4347 8672
rect 1715 8192 2035 8193
rect 1715 8128 1723 8192
rect 1787 8128 1803 8192
rect 1867 8128 1883 8192
rect 1947 8128 1963 8192
rect 2027 8128 2035 8192
rect 1715 8127 2035 8128
rect 3256 8192 3576 8193
rect 3256 8128 3264 8192
rect 3328 8128 3344 8192
rect 3408 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3576 8192
rect 3256 8127 3576 8128
rect 4798 8192 5118 8193
rect 4798 8128 4806 8192
rect 4870 8128 4886 8192
rect 4950 8128 4966 8192
rect 5030 8128 5046 8192
rect 5110 8128 5118 8192
rect 4798 8127 5118 8128
rect 2485 7648 2805 7649
rect 2485 7584 2493 7648
rect 2557 7584 2573 7648
rect 2637 7584 2653 7648
rect 2717 7584 2733 7648
rect 2797 7584 2805 7648
rect 2485 7583 2805 7584
rect 4027 7648 4347 7649
rect 4027 7584 4035 7648
rect 4099 7584 4115 7648
rect 4179 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4347 7648
rect 4027 7583 4347 7584
rect 1715 7104 2035 7105
rect 1715 7040 1723 7104
rect 1787 7040 1803 7104
rect 1867 7040 1883 7104
rect 1947 7040 1963 7104
rect 2027 7040 2035 7104
rect 1715 7039 2035 7040
rect 3256 7104 3576 7105
rect 3256 7040 3264 7104
rect 3328 7040 3344 7104
rect 3408 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3576 7104
rect 3256 7039 3576 7040
rect 4798 7104 5118 7105
rect 4798 7040 4806 7104
rect 4870 7040 4886 7104
rect 4950 7040 4966 7104
rect 5030 7040 5046 7104
rect 5110 7040 5118 7104
rect 4798 7039 5118 7040
rect 2485 6560 2805 6561
rect 2485 6496 2493 6560
rect 2557 6496 2573 6560
rect 2637 6496 2653 6560
rect 2717 6496 2733 6560
rect 2797 6496 2805 6560
rect 2485 6495 2805 6496
rect 4027 6560 4347 6561
rect 4027 6496 4035 6560
rect 4099 6496 4115 6560
rect 4179 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4347 6560
rect 4027 6495 4347 6496
rect 1715 6016 2035 6017
rect 1715 5952 1723 6016
rect 1787 5952 1803 6016
rect 1867 5952 1883 6016
rect 1947 5952 1963 6016
rect 2027 5952 2035 6016
rect 1715 5951 2035 5952
rect 3256 6016 3576 6017
rect 3256 5952 3264 6016
rect 3328 5952 3344 6016
rect 3408 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3576 6016
rect 3256 5951 3576 5952
rect 4798 6016 5118 6017
rect 4798 5952 4806 6016
rect 4870 5952 4886 6016
rect 4950 5952 4966 6016
rect 5030 5952 5046 6016
rect 5110 5952 5118 6016
rect 4798 5951 5118 5952
rect 0 5538 800 5568
rect 0 5478 1594 5538
rect 0 5448 800 5478
rect 1534 5266 1594 5478
rect 2485 5472 2805 5473
rect 2485 5408 2493 5472
rect 2557 5408 2573 5472
rect 2637 5408 2653 5472
rect 2717 5408 2733 5472
rect 2797 5408 2805 5472
rect 2485 5407 2805 5408
rect 4027 5472 4347 5473
rect 4027 5408 4035 5472
rect 4099 5408 4115 5472
rect 4179 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4347 5472
rect 4027 5407 4347 5408
rect 2957 5266 3023 5269
rect 1534 5264 3023 5266
rect 1534 5208 2962 5264
rect 3018 5208 3023 5264
rect 1534 5206 3023 5208
rect 2957 5203 3023 5206
rect 1715 4928 2035 4929
rect 1715 4864 1723 4928
rect 1787 4864 1803 4928
rect 1867 4864 1883 4928
rect 1947 4864 1963 4928
rect 2027 4864 2035 4928
rect 1715 4863 2035 4864
rect 3256 4928 3576 4929
rect 3256 4864 3264 4928
rect 3328 4864 3344 4928
rect 3408 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3576 4928
rect 3256 4863 3576 4864
rect 4798 4928 5118 4929
rect 4798 4864 4806 4928
rect 4870 4864 4886 4928
rect 4950 4864 4966 4928
rect 5030 4864 5046 4928
rect 5110 4864 5118 4928
rect 4798 4863 5118 4864
rect 5257 4858 5323 4861
rect 6033 4858 6833 4888
rect 5257 4856 6833 4858
rect 5257 4800 5262 4856
rect 5318 4800 6833 4856
rect 5257 4798 6833 4800
rect 5257 4795 5323 4798
rect 6033 4768 6833 4798
rect 2485 4384 2805 4385
rect 2485 4320 2493 4384
rect 2557 4320 2573 4384
rect 2637 4320 2653 4384
rect 2717 4320 2733 4384
rect 2797 4320 2805 4384
rect 2485 4319 2805 4320
rect 4027 4384 4347 4385
rect 4027 4320 4035 4384
rect 4099 4320 4115 4384
rect 4179 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4347 4384
rect 4027 4319 4347 4320
rect 1715 3840 2035 3841
rect 1715 3776 1723 3840
rect 1787 3776 1803 3840
rect 1867 3776 1883 3840
rect 1947 3776 1963 3840
rect 2027 3776 2035 3840
rect 1715 3775 2035 3776
rect 3256 3840 3576 3841
rect 3256 3776 3264 3840
rect 3328 3776 3344 3840
rect 3408 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3576 3840
rect 3256 3775 3576 3776
rect 4798 3840 5118 3841
rect 4798 3776 4806 3840
rect 4870 3776 4886 3840
rect 4950 3776 4966 3840
rect 5030 3776 5046 3840
rect 5110 3776 5118 3840
rect 4798 3775 5118 3776
rect 2485 3296 2805 3297
rect 2485 3232 2493 3296
rect 2557 3232 2573 3296
rect 2637 3232 2653 3296
rect 2717 3232 2733 3296
rect 2797 3232 2805 3296
rect 2485 3231 2805 3232
rect 4027 3296 4347 3297
rect 4027 3232 4035 3296
rect 4099 3232 4115 3296
rect 4179 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4347 3296
rect 4027 3231 4347 3232
rect 1715 2752 2035 2753
rect 1715 2688 1723 2752
rect 1787 2688 1803 2752
rect 1867 2688 1883 2752
rect 1947 2688 1963 2752
rect 2027 2688 2035 2752
rect 1715 2687 2035 2688
rect 3256 2752 3576 2753
rect 3256 2688 3264 2752
rect 3328 2688 3344 2752
rect 3408 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3576 2752
rect 3256 2687 3576 2688
rect 4798 2752 5118 2753
rect 4798 2688 4806 2752
rect 4870 2688 4886 2752
rect 4950 2688 4966 2752
rect 5030 2688 5046 2752
rect 5110 2688 5118 2752
rect 4798 2687 5118 2688
rect 2485 2208 2805 2209
rect 2485 2144 2493 2208
rect 2557 2144 2573 2208
rect 2637 2144 2653 2208
rect 2717 2144 2733 2208
rect 2797 2144 2805 2208
rect 2485 2143 2805 2144
rect 4027 2208 4347 2209
rect 4027 2144 4035 2208
rect 4099 2144 4115 2208
rect 4179 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4347 2208
rect 4027 2143 4347 2144
<< via3 >>
rect 2493 8732 2557 8736
rect 2493 8676 2497 8732
rect 2497 8676 2553 8732
rect 2553 8676 2557 8732
rect 2493 8672 2557 8676
rect 2573 8732 2637 8736
rect 2573 8676 2577 8732
rect 2577 8676 2633 8732
rect 2633 8676 2637 8732
rect 2573 8672 2637 8676
rect 2653 8732 2717 8736
rect 2653 8676 2657 8732
rect 2657 8676 2713 8732
rect 2713 8676 2717 8732
rect 2653 8672 2717 8676
rect 2733 8732 2797 8736
rect 2733 8676 2737 8732
rect 2737 8676 2793 8732
rect 2793 8676 2797 8732
rect 2733 8672 2797 8676
rect 4035 8732 4099 8736
rect 4035 8676 4039 8732
rect 4039 8676 4095 8732
rect 4095 8676 4099 8732
rect 4035 8672 4099 8676
rect 4115 8732 4179 8736
rect 4115 8676 4119 8732
rect 4119 8676 4175 8732
rect 4175 8676 4179 8732
rect 4115 8672 4179 8676
rect 4195 8732 4259 8736
rect 4195 8676 4199 8732
rect 4199 8676 4255 8732
rect 4255 8676 4259 8732
rect 4195 8672 4259 8676
rect 4275 8732 4339 8736
rect 4275 8676 4279 8732
rect 4279 8676 4335 8732
rect 4335 8676 4339 8732
rect 4275 8672 4339 8676
rect 1723 8188 1787 8192
rect 1723 8132 1727 8188
rect 1727 8132 1783 8188
rect 1783 8132 1787 8188
rect 1723 8128 1787 8132
rect 1803 8188 1867 8192
rect 1803 8132 1807 8188
rect 1807 8132 1863 8188
rect 1863 8132 1867 8188
rect 1803 8128 1867 8132
rect 1883 8188 1947 8192
rect 1883 8132 1887 8188
rect 1887 8132 1943 8188
rect 1943 8132 1947 8188
rect 1883 8128 1947 8132
rect 1963 8188 2027 8192
rect 1963 8132 1967 8188
rect 1967 8132 2023 8188
rect 2023 8132 2027 8188
rect 1963 8128 2027 8132
rect 3264 8188 3328 8192
rect 3264 8132 3268 8188
rect 3268 8132 3324 8188
rect 3324 8132 3328 8188
rect 3264 8128 3328 8132
rect 3344 8188 3408 8192
rect 3344 8132 3348 8188
rect 3348 8132 3404 8188
rect 3404 8132 3408 8188
rect 3344 8128 3408 8132
rect 3424 8188 3488 8192
rect 3424 8132 3428 8188
rect 3428 8132 3484 8188
rect 3484 8132 3488 8188
rect 3424 8128 3488 8132
rect 3504 8188 3568 8192
rect 3504 8132 3508 8188
rect 3508 8132 3564 8188
rect 3564 8132 3568 8188
rect 3504 8128 3568 8132
rect 4806 8188 4870 8192
rect 4806 8132 4810 8188
rect 4810 8132 4866 8188
rect 4866 8132 4870 8188
rect 4806 8128 4870 8132
rect 4886 8188 4950 8192
rect 4886 8132 4890 8188
rect 4890 8132 4946 8188
rect 4946 8132 4950 8188
rect 4886 8128 4950 8132
rect 4966 8188 5030 8192
rect 4966 8132 4970 8188
rect 4970 8132 5026 8188
rect 5026 8132 5030 8188
rect 4966 8128 5030 8132
rect 5046 8188 5110 8192
rect 5046 8132 5050 8188
rect 5050 8132 5106 8188
rect 5106 8132 5110 8188
rect 5046 8128 5110 8132
rect 2493 7644 2557 7648
rect 2493 7588 2497 7644
rect 2497 7588 2553 7644
rect 2553 7588 2557 7644
rect 2493 7584 2557 7588
rect 2573 7644 2637 7648
rect 2573 7588 2577 7644
rect 2577 7588 2633 7644
rect 2633 7588 2637 7644
rect 2573 7584 2637 7588
rect 2653 7644 2717 7648
rect 2653 7588 2657 7644
rect 2657 7588 2713 7644
rect 2713 7588 2717 7644
rect 2653 7584 2717 7588
rect 2733 7644 2797 7648
rect 2733 7588 2737 7644
rect 2737 7588 2793 7644
rect 2793 7588 2797 7644
rect 2733 7584 2797 7588
rect 4035 7644 4099 7648
rect 4035 7588 4039 7644
rect 4039 7588 4095 7644
rect 4095 7588 4099 7644
rect 4035 7584 4099 7588
rect 4115 7644 4179 7648
rect 4115 7588 4119 7644
rect 4119 7588 4175 7644
rect 4175 7588 4179 7644
rect 4115 7584 4179 7588
rect 4195 7644 4259 7648
rect 4195 7588 4199 7644
rect 4199 7588 4255 7644
rect 4255 7588 4259 7644
rect 4195 7584 4259 7588
rect 4275 7644 4339 7648
rect 4275 7588 4279 7644
rect 4279 7588 4335 7644
rect 4335 7588 4339 7644
rect 4275 7584 4339 7588
rect 1723 7100 1787 7104
rect 1723 7044 1727 7100
rect 1727 7044 1783 7100
rect 1783 7044 1787 7100
rect 1723 7040 1787 7044
rect 1803 7100 1867 7104
rect 1803 7044 1807 7100
rect 1807 7044 1863 7100
rect 1863 7044 1867 7100
rect 1803 7040 1867 7044
rect 1883 7100 1947 7104
rect 1883 7044 1887 7100
rect 1887 7044 1943 7100
rect 1943 7044 1947 7100
rect 1883 7040 1947 7044
rect 1963 7100 2027 7104
rect 1963 7044 1967 7100
rect 1967 7044 2023 7100
rect 2023 7044 2027 7100
rect 1963 7040 2027 7044
rect 3264 7100 3328 7104
rect 3264 7044 3268 7100
rect 3268 7044 3324 7100
rect 3324 7044 3328 7100
rect 3264 7040 3328 7044
rect 3344 7100 3408 7104
rect 3344 7044 3348 7100
rect 3348 7044 3404 7100
rect 3404 7044 3408 7100
rect 3344 7040 3408 7044
rect 3424 7100 3488 7104
rect 3424 7044 3428 7100
rect 3428 7044 3484 7100
rect 3484 7044 3488 7100
rect 3424 7040 3488 7044
rect 3504 7100 3568 7104
rect 3504 7044 3508 7100
rect 3508 7044 3564 7100
rect 3564 7044 3568 7100
rect 3504 7040 3568 7044
rect 4806 7100 4870 7104
rect 4806 7044 4810 7100
rect 4810 7044 4866 7100
rect 4866 7044 4870 7100
rect 4806 7040 4870 7044
rect 4886 7100 4950 7104
rect 4886 7044 4890 7100
rect 4890 7044 4946 7100
rect 4946 7044 4950 7100
rect 4886 7040 4950 7044
rect 4966 7100 5030 7104
rect 4966 7044 4970 7100
rect 4970 7044 5026 7100
rect 5026 7044 5030 7100
rect 4966 7040 5030 7044
rect 5046 7100 5110 7104
rect 5046 7044 5050 7100
rect 5050 7044 5106 7100
rect 5106 7044 5110 7100
rect 5046 7040 5110 7044
rect 2493 6556 2557 6560
rect 2493 6500 2497 6556
rect 2497 6500 2553 6556
rect 2553 6500 2557 6556
rect 2493 6496 2557 6500
rect 2573 6556 2637 6560
rect 2573 6500 2577 6556
rect 2577 6500 2633 6556
rect 2633 6500 2637 6556
rect 2573 6496 2637 6500
rect 2653 6556 2717 6560
rect 2653 6500 2657 6556
rect 2657 6500 2713 6556
rect 2713 6500 2717 6556
rect 2653 6496 2717 6500
rect 2733 6556 2797 6560
rect 2733 6500 2737 6556
rect 2737 6500 2793 6556
rect 2793 6500 2797 6556
rect 2733 6496 2797 6500
rect 4035 6556 4099 6560
rect 4035 6500 4039 6556
rect 4039 6500 4095 6556
rect 4095 6500 4099 6556
rect 4035 6496 4099 6500
rect 4115 6556 4179 6560
rect 4115 6500 4119 6556
rect 4119 6500 4175 6556
rect 4175 6500 4179 6556
rect 4115 6496 4179 6500
rect 4195 6556 4259 6560
rect 4195 6500 4199 6556
rect 4199 6500 4255 6556
rect 4255 6500 4259 6556
rect 4195 6496 4259 6500
rect 4275 6556 4339 6560
rect 4275 6500 4279 6556
rect 4279 6500 4335 6556
rect 4335 6500 4339 6556
rect 4275 6496 4339 6500
rect 1723 6012 1787 6016
rect 1723 5956 1727 6012
rect 1727 5956 1783 6012
rect 1783 5956 1787 6012
rect 1723 5952 1787 5956
rect 1803 6012 1867 6016
rect 1803 5956 1807 6012
rect 1807 5956 1863 6012
rect 1863 5956 1867 6012
rect 1803 5952 1867 5956
rect 1883 6012 1947 6016
rect 1883 5956 1887 6012
rect 1887 5956 1943 6012
rect 1943 5956 1947 6012
rect 1883 5952 1947 5956
rect 1963 6012 2027 6016
rect 1963 5956 1967 6012
rect 1967 5956 2023 6012
rect 2023 5956 2027 6012
rect 1963 5952 2027 5956
rect 3264 6012 3328 6016
rect 3264 5956 3268 6012
rect 3268 5956 3324 6012
rect 3324 5956 3328 6012
rect 3264 5952 3328 5956
rect 3344 6012 3408 6016
rect 3344 5956 3348 6012
rect 3348 5956 3404 6012
rect 3404 5956 3408 6012
rect 3344 5952 3408 5956
rect 3424 6012 3488 6016
rect 3424 5956 3428 6012
rect 3428 5956 3484 6012
rect 3484 5956 3488 6012
rect 3424 5952 3488 5956
rect 3504 6012 3568 6016
rect 3504 5956 3508 6012
rect 3508 5956 3564 6012
rect 3564 5956 3568 6012
rect 3504 5952 3568 5956
rect 4806 6012 4870 6016
rect 4806 5956 4810 6012
rect 4810 5956 4866 6012
rect 4866 5956 4870 6012
rect 4806 5952 4870 5956
rect 4886 6012 4950 6016
rect 4886 5956 4890 6012
rect 4890 5956 4946 6012
rect 4946 5956 4950 6012
rect 4886 5952 4950 5956
rect 4966 6012 5030 6016
rect 4966 5956 4970 6012
rect 4970 5956 5026 6012
rect 5026 5956 5030 6012
rect 4966 5952 5030 5956
rect 5046 6012 5110 6016
rect 5046 5956 5050 6012
rect 5050 5956 5106 6012
rect 5106 5956 5110 6012
rect 5046 5952 5110 5956
rect 2493 5468 2557 5472
rect 2493 5412 2497 5468
rect 2497 5412 2553 5468
rect 2553 5412 2557 5468
rect 2493 5408 2557 5412
rect 2573 5468 2637 5472
rect 2573 5412 2577 5468
rect 2577 5412 2633 5468
rect 2633 5412 2637 5468
rect 2573 5408 2637 5412
rect 2653 5468 2717 5472
rect 2653 5412 2657 5468
rect 2657 5412 2713 5468
rect 2713 5412 2717 5468
rect 2653 5408 2717 5412
rect 2733 5468 2797 5472
rect 2733 5412 2737 5468
rect 2737 5412 2793 5468
rect 2793 5412 2797 5468
rect 2733 5408 2797 5412
rect 4035 5468 4099 5472
rect 4035 5412 4039 5468
rect 4039 5412 4095 5468
rect 4095 5412 4099 5468
rect 4035 5408 4099 5412
rect 4115 5468 4179 5472
rect 4115 5412 4119 5468
rect 4119 5412 4175 5468
rect 4175 5412 4179 5468
rect 4115 5408 4179 5412
rect 4195 5468 4259 5472
rect 4195 5412 4199 5468
rect 4199 5412 4255 5468
rect 4255 5412 4259 5468
rect 4195 5408 4259 5412
rect 4275 5468 4339 5472
rect 4275 5412 4279 5468
rect 4279 5412 4335 5468
rect 4335 5412 4339 5468
rect 4275 5408 4339 5412
rect 1723 4924 1787 4928
rect 1723 4868 1727 4924
rect 1727 4868 1783 4924
rect 1783 4868 1787 4924
rect 1723 4864 1787 4868
rect 1803 4924 1867 4928
rect 1803 4868 1807 4924
rect 1807 4868 1863 4924
rect 1863 4868 1867 4924
rect 1803 4864 1867 4868
rect 1883 4924 1947 4928
rect 1883 4868 1887 4924
rect 1887 4868 1943 4924
rect 1943 4868 1947 4924
rect 1883 4864 1947 4868
rect 1963 4924 2027 4928
rect 1963 4868 1967 4924
rect 1967 4868 2023 4924
rect 2023 4868 2027 4924
rect 1963 4864 2027 4868
rect 3264 4924 3328 4928
rect 3264 4868 3268 4924
rect 3268 4868 3324 4924
rect 3324 4868 3328 4924
rect 3264 4864 3328 4868
rect 3344 4924 3408 4928
rect 3344 4868 3348 4924
rect 3348 4868 3404 4924
rect 3404 4868 3408 4924
rect 3344 4864 3408 4868
rect 3424 4924 3488 4928
rect 3424 4868 3428 4924
rect 3428 4868 3484 4924
rect 3484 4868 3488 4924
rect 3424 4864 3488 4868
rect 3504 4924 3568 4928
rect 3504 4868 3508 4924
rect 3508 4868 3564 4924
rect 3564 4868 3568 4924
rect 3504 4864 3568 4868
rect 4806 4924 4870 4928
rect 4806 4868 4810 4924
rect 4810 4868 4866 4924
rect 4866 4868 4870 4924
rect 4806 4864 4870 4868
rect 4886 4924 4950 4928
rect 4886 4868 4890 4924
rect 4890 4868 4946 4924
rect 4946 4868 4950 4924
rect 4886 4864 4950 4868
rect 4966 4924 5030 4928
rect 4966 4868 4970 4924
rect 4970 4868 5026 4924
rect 5026 4868 5030 4924
rect 4966 4864 5030 4868
rect 5046 4924 5110 4928
rect 5046 4868 5050 4924
rect 5050 4868 5106 4924
rect 5106 4868 5110 4924
rect 5046 4864 5110 4868
rect 2493 4380 2557 4384
rect 2493 4324 2497 4380
rect 2497 4324 2553 4380
rect 2553 4324 2557 4380
rect 2493 4320 2557 4324
rect 2573 4380 2637 4384
rect 2573 4324 2577 4380
rect 2577 4324 2633 4380
rect 2633 4324 2637 4380
rect 2573 4320 2637 4324
rect 2653 4380 2717 4384
rect 2653 4324 2657 4380
rect 2657 4324 2713 4380
rect 2713 4324 2717 4380
rect 2653 4320 2717 4324
rect 2733 4380 2797 4384
rect 2733 4324 2737 4380
rect 2737 4324 2793 4380
rect 2793 4324 2797 4380
rect 2733 4320 2797 4324
rect 4035 4380 4099 4384
rect 4035 4324 4039 4380
rect 4039 4324 4095 4380
rect 4095 4324 4099 4380
rect 4035 4320 4099 4324
rect 4115 4380 4179 4384
rect 4115 4324 4119 4380
rect 4119 4324 4175 4380
rect 4175 4324 4179 4380
rect 4115 4320 4179 4324
rect 4195 4380 4259 4384
rect 4195 4324 4199 4380
rect 4199 4324 4255 4380
rect 4255 4324 4259 4380
rect 4195 4320 4259 4324
rect 4275 4380 4339 4384
rect 4275 4324 4279 4380
rect 4279 4324 4335 4380
rect 4335 4324 4339 4380
rect 4275 4320 4339 4324
rect 1723 3836 1787 3840
rect 1723 3780 1727 3836
rect 1727 3780 1783 3836
rect 1783 3780 1787 3836
rect 1723 3776 1787 3780
rect 1803 3836 1867 3840
rect 1803 3780 1807 3836
rect 1807 3780 1863 3836
rect 1863 3780 1867 3836
rect 1803 3776 1867 3780
rect 1883 3836 1947 3840
rect 1883 3780 1887 3836
rect 1887 3780 1943 3836
rect 1943 3780 1947 3836
rect 1883 3776 1947 3780
rect 1963 3836 2027 3840
rect 1963 3780 1967 3836
rect 1967 3780 2023 3836
rect 2023 3780 2027 3836
rect 1963 3776 2027 3780
rect 3264 3836 3328 3840
rect 3264 3780 3268 3836
rect 3268 3780 3324 3836
rect 3324 3780 3328 3836
rect 3264 3776 3328 3780
rect 3344 3836 3408 3840
rect 3344 3780 3348 3836
rect 3348 3780 3404 3836
rect 3404 3780 3408 3836
rect 3344 3776 3408 3780
rect 3424 3836 3488 3840
rect 3424 3780 3428 3836
rect 3428 3780 3484 3836
rect 3484 3780 3488 3836
rect 3424 3776 3488 3780
rect 3504 3836 3568 3840
rect 3504 3780 3508 3836
rect 3508 3780 3564 3836
rect 3564 3780 3568 3836
rect 3504 3776 3568 3780
rect 4806 3836 4870 3840
rect 4806 3780 4810 3836
rect 4810 3780 4866 3836
rect 4866 3780 4870 3836
rect 4806 3776 4870 3780
rect 4886 3836 4950 3840
rect 4886 3780 4890 3836
rect 4890 3780 4946 3836
rect 4946 3780 4950 3836
rect 4886 3776 4950 3780
rect 4966 3836 5030 3840
rect 4966 3780 4970 3836
rect 4970 3780 5026 3836
rect 5026 3780 5030 3836
rect 4966 3776 5030 3780
rect 5046 3836 5110 3840
rect 5046 3780 5050 3836
rect 5050 3780 5106 3836
rect 5106 3780 5110 3836
rect 5046 3776 5110 3780
rect 2493 3292 2557 3296
rect 2493 3236 2497 3292
rect 2497 3236 2553 3292
rect 2553 3236 2557 3292
rect 2493 3232 2557 3236
rect 2573 3292 2637 3296
rect 2573 3236 2577 3292
rect 2577 3236 2633 3292
rect 2633 3236 2637 3292
rect 2573 3232 2637 3236
rect 2653 3292 2717 3296
rect 2653 3236 2657 3292
rect 2657 3236 2713 3292
rect 2713 3236 2717 3292
rect 2653 3232 2717 3236
rect 2733 3292 2797 3296
rect 2733 3236 2737 3292
rect 2737 3236 2793 3292
rect 2793 3236 2797 3292
rect 2733 3232 2797 3236
rect 4035 3292 4099 3296
rect 4035 3236 4039 3292
rect 4039 3236 4095 3292
rect 4095 3236 4099 3292
rect 4035 3232 4099 3236
rect 4115 3292 4179 3296
rect 4115 3236 4119 3292
rect 4119 3236 4175 3292
rect 4175 3236 4179 3292
rect 4115 3232 4179 3236
rect 4195 3292 4259 3296
rect 4195 3236 4199 3292
rect 4199 3236 4255 3292
rect 4255 3236 4259 3292
rect 4195 3232 4259 3236
rect 4275 3292 4339 3296
rect 4275 3236 4279 3292
rect 4279 3236 4335 3292
rect 4335 3236 4339 3292
rect 4275 3232 4339 3236
rect 1723 2748 1787 2752
rect 1723 2692 1727 2748
rect 1727 2692 1783 2748
rect 1783 2692 1787 2748
rect 1723 2688 1787 2692
rect 1803 2748 1867 2752
rect 1803 2692 1807 2748
rect 1807 2692 1863 2748
rect 1863 2692 1867 2748
rect 1803 2688 1867 2692
rect 1883 2748 1947 2752
rect 1883 2692 1887 2748
rect 1887 2692 1943 2748
rect 1943 2692 1947 2748
rect 1883 2688 1947 2692
rect 1963 2748 2027 2752
rect 1963 2692 1967 2748
rect 1967 2692 2023 2748
rect 2023 2692 2027 2748
rect 1963 2688 2027 2692
rect 3264 2748 3328 2752
rect 3264 2692 3268 2748
rect 3268 2692 3324 2748
rect 3324 2692 3328 2748
rect 3264 2688 3328 2692
rect 3344 2748 3408 2752
rect 3344 2692 3348 2748
rect 3348 2692 3404 2748
rect 3404 2692 3408 2748
rect 3344 2688 3408 2692
rect 3424 2748 3488 2752
rect 3424 2692 3428 2748
rect 3428 2692 3484 2748
rect 3484 2692 3488 2748
rect 3424 2688 3488 2692
rect 3504 2748 3568 2752
rect 3504 2692 3508 2748
rect 3508 2692 3564 2748
rect 3564 2692 3568 2748
rect 3504 2688 3568 2692
rect 4806 2748 4870 2752
rect 4806 2692 4810 2748
rect 4810 2692 4866 2748
rect 4866 2692 4870 2748
rect 4806 2688 4870 2692
rect 4886 2748 4950 2752
rect 4886 2692 4890 2748
rect 4890 2692 4946 2748
rect 4946 2692 4950 2748
rect 4886 2688 4950 2692
rect 4966 2748 5030 2752
rect 4966 2692 4970 2748
rect 4970 2692 5026 2748
rect 5026 2692 5030 2748
rect 4966 2688 5030 2692
rect 5046 2748 5110 2752
rect 5046 2692 5050 2748
rect 5050 2692 5106 2748
rect 5106 2692 5110 2748
rect 5046 2688 5110 2692
rect 2493 2204 2557 2208
rect 2493 2148 2497 2204
rect 2497 2148 2553 2204
rect 2553 2148 2557 2204
rect 2493 2144 2557 2148
rect 2573 2204 2637 2208
rect 2573 2148 2577 2204
rect 2577 2148 2633 2204
rect 2633 2148 2637 2204
rect 2573 2144 2637 2148
rect 2653 2204 2717 2208
rect 2653 2148 2657 2204
rect 2657 2148 2713 2204
rect 2713 2148 2717 2204
rect 2653 2144 2717 2148
rect 2733 2204 2797 2208
rect 2733 2148 2737 2204
rect 2737 2148 2793 2204
rect 2793 2148 2797 2204
rect 2733 2144 2797 2148
rect 4035 2204 4099 2208
rect 4035 2148 4039 2204
rect 4039 2148 4095 2204
rect 4095 2148 4099 2204
rect 4035 2144 4099 2148
rect 4115 2204 4179 2208
rect 4115 2148 4119 2204
rect 4119 2148 4175 2204
rect 4175 2148 4179 2204
rect 4115 2144 4179 2148
rect 4195 2204 4259 2208
rect 4195 2148 4199 2204
rect 4199 2148 4255 2204
rect 4255 2148 4259 2204
rect 4195 2144 4259 2148
rect 4275 2204 4339 2208
rect 4275 2148 4279 2204
rect 4279 2148 4335 2204
rect 4335 2148 4339 2204
rect 4275 2144 4339 2148
<< metal4 >>
rect 1715 8192 2035 8752
rect 1715 8128 1723 8192
rect 1787 8128 1803 8192
rect 1867 8128 1883 8192
rect 1947 8128 1963 8192
rect 2027 8128 2035 8192
rect 1715 7767 2035 8128
rect 1715 7531 1757 7767
rect 1993 7531 2035 7767
rect 1715 7104 2035 7531
rect 1715 7040 1723 7104
rect 1787 7040 1803 7104
rect 1867 7040 1883 7104
rect 1947 7040 1963 7104
rect 2027 7040 2035 7104
rect 1715 6016 2035 7040
rect 1715 5952 1723 6016
rect 1787 5952 1803 6016
rect 1867 5952 1883 6016
rect 1947 5952 1963 6016
rect 2027 5952 2035 6016
rect 1715 5558 2035 5952
rect 1715 5322 1757 5558
rect 1993 5322 2035 5558
rect 1715 4928 2035 5322
rect 1715 4864 1723 4928
rect 1787 4864 1803 4928
rect 1867 4864 1883 4928
rect 1947 4864 1963 4928
rect 2027 4864 2035 4928
rect 1715 3840 2035 4864
rect 1715 3776 1723 3840
rect 1787 3776 1803 3840
rect 1867 3776 1883 3840
rect 1947 3776 1963 3840
rect 2027 3776 2035 3840
rect 1715 3350 2035 3776
rect 1715 3114 1757 3350
rect 1993 3114 2035 3350
rect 1715 2752 2035 3114
rect 1715 2688 1723 2752
rect 1787 2688 1803 2752
rect 1867 2688 1883 2752
rect 1947 2688 1963 2752
rect 2027 2688 2035 2752
rect 1715 2128 2035 2688
rect 2485 8736 2805 8752
rect 2485 8672 2493 8736
rect 2557 8672 2573 8736
rect 2637 8672 2653 8736
rect 2717 8672 2733 8736
rect 2797 8672 2805 8736
rect 2485 7648 2805 8672
rect 2485 7584 2493 7648
rect 2557 7584 2573 7648
rect 2637 7584 2653 7648
rect 2717 7584 2733 7648
rect 2797 7584 2805 7648
rect 2485 6663 2805 7584
rect 2485 6560 2527 6663
rect 2763 6560 2805 6663
rect 2485 6496 2493 6560
rect 2797 6496 2805 6560
rect 2485 6427 2527 6496
rect 2763 6427 2805 6496
rect 2485 5472 2805 6427
rect 2485 5408 2493 5472
rect 2557 5408 2573 5472
rect 2637 5408 2653 5472
rect 2717 5408 2733 5472
rect 2797 5408 2805 5472
rect 2485 4454 2805 5408
rect 2485 4384 2527 4454
rect 2763 4384 2805 4454
rect 2485 4320 2493 4384
rect 2797 4320 2805 4384
rect 2485 4218 2527 4320
rect 2763 4218 2805 4320
rect 2485 3296 2805 4218
rect 2485 3232 2493 3296
rect 2557 3232 2573 3296
rect 2637 3232 2653 3296
rect 2717 3232 2733 3296
rect 2797 3232 2805 3296
rect 2485 2208 2805 3232
rect 2485 2144 2493 2208
rect 2557 2144 2573 2208
rect 2637 2144 2653 2208
rect 2717 2144 2733 2208
rect 2797 2144 2805 2208
rect 2485 2128 2805 2144
rect 3256 8192 3576 8752
rect 3256 8128 3264 8192
rect 3328 8128 3344 8192
rect 3408 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3576 8192
rect 3256 7767 3576 8128
rect 3256 7531 3298 7767
rect 3534 7531 3576 7767
rect 3256 7104 3576 7531
rect 3256 7040 3264 7104
rect 3328 7040 3344 7104
rect 3408 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3576 7104
rect 3256 6016 3576 7040
rect 3256 5952 3264 6016
rect 3328 5952 3344 6016
rect 3408 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3576 6016
rect 3256 5558 3576 5952
rect 3256 5322 3298 5558
rect 3534 5322 3576 5558
rect 3256 4928 3576 5322
rect 3256 4864 3264 4928
rect 3328 4864 3344 4928
rect 3408 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3576 4928
rect 3256 3840 3576 4864
rect 3256 3776 3264 3840
rect 3328 3776 3344 3840
rect 3408 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3576 3840
rect 3256 3350 3576 3776
rect 3256 3114 3298 3350
rect 3534 3114 3576 3350
rect 3256 2752 3576 3114
rect 3256 2688 3264 2752
rect 3328 2688 3344 2752
rect 3408 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3576 2752
rect 3256 2128 3576 2688
rect 4027 8736 4347 8752
rect 4027 8672 4035 8736
rect 4099 8672 4115 8736
rect 4179 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4347 8736
rect 4027 7648 4347 8672
rect 4027 7584 4035 7648
rect 4099 7584 4115 7648
rect 4179 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4347 7648
rect 4027 6663 4347 7584
rect 4027 6560 4069 6663
rect 4305 6560 4347 6663
rect 4027 6496 4035 6560
rect 4339 6496 4347 6560
rect 4027 6427 4069 6496
rect 4305 6427 4347 6496
rect 4027 5472 4347 6427
rect 4027 5408 4035 5472
rect 4099 5408 4115 5472
rect 4179 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4347 5472
rect 4027 4454 4347 5408
rect 4027 4384 4069 4454
rect 4305 4384 4347 4454
rect 4027 4320 4035 4384
rect 4339 4320 4347 4384
rect 4027 4218 4069 4320
rect 4305 4218 4347 4320
rect 4027 3296 4347 4218
rect 4027 3232 4035 3296
rect 4099 3232 4115 3296
rect 4179 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4347 3296
rect 4027 2208 4347 3232
rect 4027 2144 4035 2208
rect 4099 2144 4115 2208
rect 4179 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4347 2208
rect 4027 2128 4347 2144
rect 4798 8192 5118 8752
rect 4798 8128 4806 8192
rect 4870 8128 4886 8192
rect 4950 8128 4966 8192
rect 5030 8128 5046 8192
rect 5110 8128 5118 8192
rect 4798 7767 5118 8128
rect 4798 7531 4840 7767
rect 5076 7531 5118 7767
rect 4798 7104 5118 7531
rect 4798 7040 4806 7104
rect 4870 7040 4886 7104
rect 4950 7040 4966 7104
rect 5030 7040 5046 7104
rect 5110 7040 5118 7104
rect 4798 6016 5118 7040
rect 4798 5952 4806 6016
rect 4870 5952 4886 6016
rect 4950 5952 4966 6016
rect 5030 5952 5046 6016
rect 5110 5952 5118 6016
rect 4798 5558 5118 5952
rect 4798 5322 4840 5558
rect 5076 5322 5118 5558
rect 4798 4928 5118 5322
rect 4798 4864 4806 4928
rect 4870 4864 4886 4928
rect 4950 4864 4966 4928
rect 5030 4864 5046 4928
rect 5110 4864 5118 4928
rect 4798 3840 5118 4864
rect 4798 3776 4806 3840
rect 4870 3776 4886 3840
rect 4950 3776 4966 3840
rect 5030 3776 5046 3840
rect 5110 3776 5118 3840
rect 4798 3350 5118 3776
rect 4798 3114 4840 3350
rect 5076 3114 5118 3350
rect 4798 2752 5118 3114
rect 4798 2688 4806 2752
rect 4870 2688 4886 2752
rect 4950 2688 4966 2752
rect 5030 2688 5046 2752
rect 5110 2688 5118 2752
rect 4798 2128 5118 2688
<< via4 >>
rect 1757 7531 1993 7767
rect 1757 5322 1993 5558
rect 1757 3114 1993 3350
rect 2527 6560 2763 6663
rect 2527 6496 2557 6560
rect 2557 6496 2573 6560
rect 2573 6496 2637 6560
rect 2637 6496 2653 6560
rect 2653 6496 2717 6560
rect 2717 6496 2733 6560
rect 2733 6496 2763 6560
rect 2527 6427 2763 6496
rect 2527 4384 2763 4454
rect 2527 4320 2557 4384
rect 2557 4320 2573 4384
rect 2573 4320 2637 4384
rect 2637 4320 2653 4384
rect 2653 4320 2717 4384
rect 2717 4320 2733 4384
rect 2733 4320 2763 4384
rect 2527 4218 2763 4320
rect 3298 7531 3534 7767
rect 3298 5322 3534 5558
rect 3298 3114 3534 3350
rect 4069 6560 4305 6663
rect 4069 6496 4099 6560
rect 4099 6496 4115 6560
rect 4115 6496 4179 6560
rect 4179 6496 4195 6560
rect 4195 6496 4259 6560
rect 4259 6496 4275 6560
rect 4275 6496 4305 6560
rect 4069 6427 4305 6496
rect 4069 4384 4305 4454
rect 4069 4320 4099 4384
rect 4099 4320 4115 4384
rect 4115 4320 4179 4384
rect 4179 4320 4195 4384
rect 4195 4320 4259 4384
rect 4259 4320 4275 4384
rect 4275 4320 4305 4384
rect 4069 4218 4305 4320
rect 4840 7531 5076 7767
rect 4840 5322 5076 5558
rect 4840 3114 5076 3350
<< metal5 >>
rect 1104 7767 5704 7809
rect 1104 7531 1757 7767
rect 1993 7531 3298 7767
rect 3534 7531 4840 7767
rect 5076 7531 5704 7767
rect 1104 7489 5704 7531
rect 1104 6663 5704 6705
rect 1104 6427 2527 6663
rect 2763 6427 4069 6663
rect 4305 6427 5704 6663
rect 1104 6385 5704 6427
rect 1104 5558 5704 5601
rect 1104 5322 1757 5558
rect 1993 5322 3298 5558
rect 3534 5322 4840 5558
rect 5076 5322 5704 5558
rect 1104 5280 5704 5322
rect 1104 4454 5704 4496
rect 1104 4218 2527 4454
rect 2763 4218 4069 4454
rect 4305 4218 5704 4454
rect 1104 4176 5704 4218
rect 1104 3350 5704 3392
rect 1104 3114 1757 3350
rect 1993 3114 3298 3350
rect 3534 3114 4840 3350
rect 5076 3114 5704 3350
rect 1104 3072 5704 3114
use sky130_fd_sc_hd__decap_8  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 1748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1640615124
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1640615124
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1640615124
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29
timestamp 1640615124
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1640615124
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_39
timestamp 1640615124
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 1640615124
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1640615124
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1640615124
transform -1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1640615124
transform -1 0 5704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1640615124
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_17
timestamp 1640615124
transform 1 0 2668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1640615124
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1640615124
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform -1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1640615124
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1640615124
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_39
timestamp 1640615124
transform 1 0 4692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1640615124
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1640615124
transform -1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 2392 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1640615124
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1640615124
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1640615124
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13_
timestamp 1640615124
transform -1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 2024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_23
timestamp 1640615124
transform 1 0 3220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 3588 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_43
timestamp 1640615124
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1640615124
transform -1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1640615124
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1640615124
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _26_
timestamp 1640615124
transform -1 0 3036 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1640615124
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1640615124
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_38
timestamp 1640615124
transform 1 0 4600 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1640615124
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform -1 0 4600 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_46
timestamp 1640615124
transform 1 0 5336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1640615124
transform -1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1640615124
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1640615124
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1640615124
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1640615124
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 2024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 2944 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_5_40
timestamp 1640615124
transform 1 0 4784 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_46
timestamp 1640615124
transform 1 0 5336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1640615124
transform -1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1640615124
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1640615124
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_14
timestamp 1640615124
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1640615124
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1640615124
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1640615124
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _14_
timestamp 1640615124
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _25_
timestamp 1640615124
transform -1 0 4232 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _27_
timestamp 1640615124
transform -1 0 3312 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1640615124
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_38
timestamp 1640615124
transform 1 0 4600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1640615124
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1640615124
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640615124
transform 1 0 4600 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _23_
timestamp 1640615124
transform -1 0 4600 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1640615124
transform 1 0 5336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_43
timestamp 1640615124
transform 1 0 5060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1640615124
transform -1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1640615124
transform -1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_13
timestamp 1640615124
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1640615124
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1640615124
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1640615124
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _19_
timestamp 1640615124
transform -1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1640615124
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1640615124
transform 1 0 4048 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1640615124
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _16_
timestamp 1640615124
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk_i
timestamp 1640615124
transform -1 0 4968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_42
timestamp 1640615124
transform 1 0 4968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_46
timestamp 1640615124
transform 1 0 5336 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1640615124
transform -1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1640615124
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1640615124
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1640615124
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1640615124
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_35
timestamp 1640615124
transform 1 0 4324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_39
timestamp 1640615124
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _22_
timestamp 1640615124
transform -1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1640615124
transform -1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1640615124
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1640615124
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1640615124
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1640615124
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1640615124
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_41
timestamp 1640615124
transform 1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1640615124
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1640615124
transform -1 0 5704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_19
timestamp 1640615124
transform 1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_7
timestamp 1640615124
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1640615124
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1640615124
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp 1640615124
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_29
timestamp 1640615124
transform 1 0 3772 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_37
timestamp 1640615124
transform 1 0 4508 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1640615124
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1640615124
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_43
timestamp 1640615124
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1640615124
transform -1 0 5704 0 -1 8704
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 4176 5704 4496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 6385 5704 6705 6 VGND
port 0 nsew ground input
rlabel metal4 s 2485 2128 2805 8752 6 VGND
port 0 nsew ground input
rlabel metal4 s 4027 2128 4347 8752 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 3072 5704 3392 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 5281 5704 5601 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 7489 5704 7809 6 VPWR
port 1 nsew power input
rlabel metal4 s 1715 2128 2035 8752 6 VPWR
port 1 nsew power input
rlabel metal4 s 3256 2128 3576 8752 6 VPWR
port 1 nsew power input
rlabel metal4 s 4798 2128 5118 8752 6 VPWR
port 1 nsew power input
rlabel metal3 s 0 5448 800 5568 6 clk_i
port 2 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 out_o[0]
port 3 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 out_o[1]
port 4 nsew signal tristate
rlabel metal2 s 662 10177 718 10977 6 out_o[2]
port 5 nsew signal tristate
rlabel metal2 s 6458 10177 6514 10977 6 out_o[3]
port 6 nsew signal tristate
rlabel metal3 s 6033 4768 6833 4888 6 reset_i
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 6833 10977
<< end >>
